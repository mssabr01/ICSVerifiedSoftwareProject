/*
 * Copyright 2017, Data61
 * Commonwealth Scientific and Industrial Research Organisation (CSIRO)
 * ABN 41 687 119 230.
 *
 * This software may be distributed and modified according to the terms of
 * the BSD 2-Clause license. Note that NO WARRANTY is provided.
 * See "LICENSE_BSD2.txt" for details.
 *
 * @TAG(DATA61_BSD)
 */

arch x86_64

objects {
conn1.conn6_ep = ep
conn2.conn5_ep = ep
conn3.conn7_ep = ep
conn4.conn8_ep = ep
crypto_6_0_control_9_tcb = tcb (addr: 0x53dc00,ip: 0x407931,sp: 0x52f000,elf: crypto_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [1],fault_ep: 0x00000002)
crypto_6_0_fault_handler_15_0000_tcb = tcb (addr: 0x543c00,ip: 0x407931,sp: 0x53b000,elf: crypto_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [5])
crypto_6_crypto_iface_12_0000_tcb = tcb (addr: 0x540c00,ip: 0x407931,sp: 0x535000,elf: crypto_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [3],fault_ep: 0x00000004)
crypto_cnode = cnode (4 bits)
crypto_fault_ep = ep
crypto_frame__camkes_ipc_buffer_crypto_0_control = frame (4k)
crypto_frame__camkes_ipc_buffer_crypto_0_fault_handler_0000 = frame (4k)
crypto_frame__camkes_ipc_buffer_crypto_crypto_iface_0000 = frame (4k)
crypto_group_bin_pd = pml4
crypto_interface_init_ep = ep
crypto_post_init_ep = ep
crypto_pre_init_ep = ep
frame_crypto_group_bin_0000 = frame (4k)
frame_crypto_group_bin_0001 = frame (4k)
frame_crypto_group_bin_0002 = frame (4k)
frame_crypto_group_bin_0003 = frame (4k)
frame_crypto_group_bin_0004 = frame (4k)
frame_crypto_group_bin_0005 = frame (4k)
frame_crypto_group_bin_0006 = frame (4k)
frame_crypto_group_bin_0007 = frame (4k)
frame_crypto_group_bin_0008 = frame (4k)
frame_crypto_group_bin_0009 = frame (4k)
frame_crypto_group_bin_0010 = frame (4k)
frame_crypto_group_bin_0011 = frame (4k)
frame_crypto_group_bin_0012 = frame (4k)
frame_crypto_group_bin_0013 = frame (4k)
frame_crypto_group_bin_0014 = frame (4k)
frame_crypto_group_bin_0015 = frame (4k)
frame_crypto_group_bin_0016 = frame (4k)
frame_crypto_group_bin_0017 = frame (4k)
frame_crypto_group_bin_0018 = frame (4k)
frame_crypto_group_bin_0019 = frame (4k)
frame_crypto_group_bin_0020 = frame (4k)
frame_crypto_group_bin_0021 = frame (4k)
frame_crypto_group_bin_0022 = frame (4k)
frame_crypto_group_bin_0023 = frame (4k)
frame_crypto_group_bin_0024 = frame (4k)
frame_crypto_group_bin_0025 = frame (4k)
frame_crypto_group_bin_0026 = frame (4k)
frame_crypto_group_bin_0027 = frame (4k)
frame_crypto_group_bin_0028 = frame (4k)
frame_crypto_group_bin_0029 = frame (4k)
frame_crypto_group_bin_0030 = frame (4k)
frame_crypto_group_bin_0031 = frame (4k)
frame_crypto_group_bin_0032 = frame (4k)
frame_crypto_group_bin_0035 = frame (4k)
frame_crypto_group_bin_0037 = frame (4k)
frame_crypto_group_bin_0038 = frame (4k)
frame_crypto_group_bin_0039 = frame (4k)
frame_crypto_group_bin_0041 = frame (4k)
frame_crypto_group_bin_0042 = frame (4k)
frame_crypto_group_bin_0043 = frame (4k)
frame_crypto_group_bin_0044 = frame (4k)
frame_crypto_group_bin_0045 = frame (4k)
frame_crypto_group_bin_0046 = frame (4k)
frame_crypto_group_bin_0047 = frame (4k)
frame_crypto_group_bin_0048 = frame (4k)
frame_crypto_group_bin_0049 = frame (4k)
frame_crypto_group_bin_0051 = frame (4k)
frame_crypto_group_bin_0052 = frame (4k)
frame_crypto_group_bin_0053 = frame (4k)
frame_crypto_group_bin_0054 = frame (4k)
frame_crypto_group_bin_0055 = frame (4k)
frame_crypto_group_bin_0056 = frame (4k)
frame_crypto_group_bin_0057 = frame (4k)
frame_crypto_group_bin_0058 = frame (4k)
frame_crypto_group_bin_0059 = frame (4k)
frame_crypto_group_bin_0060 = frame (4k)
frame_crypto_group_bin_0061 = frame (4k)
frame_crypto_group_bin_0062 = frame (4k)
frame_crypto_group_bin_0063 = frame (4k)
frame_crypto_group_bin_0065 = frame (4k)
frame_crypto_group_bin_0067 = frame (4k)
frame_crypto_group_bin_0068 = frame (4k)
frame_crypto_group_bin_0070 = frame (4k)
frame_crypto_group_bin_0071 = frame (4k)
frame_crypto_group_bin_0072 = frame (4k)
frame_crypto_group_bin_0073 = frame (4k)
frame_crypto_group_bin_0074 = frame (4k)
frame_crypto_group_bin_0075 = frame (4k)
frame_crypto_group_bin_0076 = frame (4k)
frame_crypto_group_bin_0077 = frame (4k)
frame_crypto_group_bin_0078 = frame (4k)
frame_crypto_group_bin_0080 = frame (4k)
frame_crypto_group_bin_0081 = frame (4k)
frame_crypto_group_bin_0083 = frame (4k)
frame_crypto_group_bin_0084 = frame (4k)
frame_crypto_group_bin_0085 = frame (4k)
frame_crypto_group_bin_0086 = frame (4k)
frame_crypto_group_bin_0087 = frame (4k)
frame_crypto_group_bin_0088 = frame (4k)
frame_crypto_group_bin_0089 = frame (4k)
frame_crypto_group_bin_0090 = frame (4k)
frame_crypto_group_bin_0091 = frame (4k)
frame_crypto_group_bin_0092 = frame (4k)
frame_crypto_group_bin_0093 = frame (4k)
frame_crypto_group_bin_0094 = frame (4k)
frame_crypto_group_bin_0095 = frame (4k)
frame_crypto_group_bin_0096 = frame (4k)
frame_crypto_group_bin_0097 = frame (4k)
frame_crypto_group_bin_0098 = frame (4k)
frame_crypto_group_bin_0099 = frame (4k)
frame_crypto_group_bin_0100 = frame (4k)
frame_crypto_group_bin_0101 = frame (4k)
frame_crypto_group_bin_0102 = frame (4k)
frame_crypto_group_bin_0104 = frame (4k)
frame_crypto_group_bin_0105 = frame (4k)
frame_crypto_group_bin_0106 = frame (4k)
frame_crypto_group_bin_0107 = frame (4k)
frame_crypto_group_bin_0108 = frame (4k)
frame_crypto_group_bin_0109 = frame (4k)
frame_crypto_group_bin_0111 = frame (4k)
frame_crypto_group_bin_0112 = frame (4k)
frame_crypto_group_bin_0114 = frame (4k)
frame_crypto_group_bin_0115 = frame (4k)
frame_crypto_group_bin_0116 = frame (4k)
frame_crypto_group_bin_0117 = frame (4k)
frame_crypto_group_bin_0118 = frame (4k)
frame_crypto_group_bin_0119 = frame (4k)
frame_crypto_group_bin_0120 = frame (4k)
frame_crypto_group_bin_0121 = frame (4k)
frame_crypto_group_bin_0122 = frame (4k)
frame_crypto_group_bin_0123 = frame (4k)
frame_crypto_group_bin_0124 = frame (4k)
frame_crypto_group_bin_0125 = frame (4k)
frame_crypto_group_bin_0126 = frame (4k)
frame_crypto_group_bin_0127 = frame (4k)
frame_crypto_group_bin_0128 = frame (4k)
frame_crypto_group_bin_0129 = frame (4k)
frame_crypto_group_bin_0130 = frame (4k)
frame_crypto_group_bin_0131 = frame (4k)
frame_crypto_group_bin_0132 = frame (4k)
frame_crypto_group_bin_0133 = frame (4k)
frame_crypto_group_bin_0134 = frame (4k)
frame_crypto_group_bin_0136 = frame (4k)
frame_crypto_group_bin_0137 = frame (4k)
frame_crypto_group_bin_0138 = frame (4k)
frame_crypto_group_bin_0139 = frame (4k)
frame_crypto_group_bin_0140 = frame (4k)
frame_crypto_group_bin_0141 = frame (4k)
frame_crypto_group_bin_0142 = frame (4k)
frame_crypto_group_bin_0143 = frame (4k)
frame_crypto_group_bin_0144 = frame (4k)
frame_crypto_group_bin_0145 = frame (4k)
frame_crypto_group_bin_0146 = frame (4k)
frame_crypto_group_bin_0147 = frame (4k)
frame_crypto_group_bin_0148 = frame (4k)
frame_crypto_group_bin_0149 = frame (4k)
frame_crypto_group_bin_0151 = frame (4k)
frame_crypto_group_bin_0152 = frame (4k)
frame_crypto_group_bin_0153 = frame (4k)
frame_crypto_group_bin_0154 = frame (4k)
frame_crypto_group_bin_0155 = frame (4k)
frame_crypto_group_bin_0156 = frame (4k)
frame_crypto_group_bin_0158 = frame (4k)
frame_crypto_group_bin_0159 = frame (4k)
frame_crypto_group_bin_0160 = frame (4k)
frame_crypto_group_bin_0161 = frame (4k)
frame_crypto_group_bin_0162 = frame (4k)
frame_crypto_group_bin_0163 = frame (4k)
frame_crypto_group_bin_0164 = frame (4k)
frame_crypto_group_bin_0165 = frame (4k)
frame_crypto_group_bin_0166 = frame (4k)
frame_crypto_group_bin_0167 = frame (4k)
frame_crypto_group_bin_0168 = frame (4k)
frame_crypto_group_bin_0169 = frame (4k)
frame_crypto_group_bin_0170 = frame (4k)
frame_crypto_group_bin_0171 = frame (4k)
frame_crypto_group_bin_0172 = frame (4k)
frame_crypto_group_bin_0174 = frame (4k)
frame_crypto_group_bin_0175 = frame (4k)
frame_crypto_group_bin_0177 = frame (4k)
frame_crypto_group_bin_0178 = frame (4k)
frame_crypto_group_bin_0179 = frame (4k)
frame_crypto_group_bin_0180 = frame (4k)
frame_crypto_group_bin_0181 = frame (4k)
frame_crypto_group_bin_0182 = frame (4k)
frame_crypto_group_bin_0184 = frame (4k)
frame_crypto_group_bin_0185 = frame (4k)
frame_crypto_group_bin_0186 = frame (4k)
frame_crypto_group_bin_0187 = frame (4k)
frame_crypto_group_bin_0188 = frame (4k)
frame_crypto_group_bin_0189 = frame (4k)
frame_crypto_group_bin_0190 = frame (4k)
frame_crypto_group_bin_0191 = frame (4k)
frame_crypto_group_bin_0192 = frame (4k)
frame_crypto_group_bin_0193 = frame (4k)
frame_crypto_group_bin_0194 = frame (4k)
frame_crypto_group_bin_0195 = frame (4k)
frame_crypto_group_bin_0196 = frame (4k)
frame_crypto_group_bin_0197 = frame (4k)
frame_crypto_group_bin_0198 = frame (4k)
frame_crypto_group_bin_0199 = frame (4k)
frame_crypto_group_bin_0200 = frame (4k)
frame_crypto_group_bin_0201 = frame (4k)
frame_crypto_group_bin_0202 = frame (4k)
frame_crypto_group_bin_0203 = frame (4k)
frame_crypto_group_bin_0204 = frame (4k)
frame_crypto_group_bin_0205 = frame (4k)
frame_crypto_group_bin_0206 = frame (4k)
frame_crypto_group_bin_0207 = frame (4k)
frame_crypto_group_bin_0208 = frame (4k)
frame_crypto_group_bin_0209 = frame (4k)
frame_crypto_group_bin_0210 = frame (4k)
frame_crypto_group_bin_0211 = frame (4k)
frame_crypto_group_bin_0212 = frame (4k)
frame_crypto_group_bin_0213 = frame (4k)
frame_crypto_group_bin_0214 = frame (4k)
frame_crypto_group_bin_0215 = frame (4k)
frame_crypto_group_bin_0216 = frame (4k)
frame_crypto_group_bin_0217 = frame (4k)
frame_crypto_group_bin_0218 = frame (4k)
frame_crypto_group_bin_0219 = frame (4k)
frame_crypto_group_bin_0221 = frame (4k)
frame_crypto_group_bin_0222 = frame (4k)
frame_crypto_group_bin_0223 = frame (4k)
frame_crypto_group_bin_0224 = frame (4k)
frame_crypto_group_bin_0225 = frame (4k)
frame_crypto_group_bin_0226 = frame (4k)
frame_crypto_group_bin_0227 = frame (4k)
frame_crypto_group_bin_0229 = frame (4k)
frame_crypto_group_bin_0230 = frame (4k)
frame_crypto_group_bin_0231 = frame (4k)
frame_crypto_group_bin_0232 = frame (4k)
frame_crypto_group_bin_0233 = frame (4k)
frame_crypto_group_bin_0234 = frame (4k)
frame_crypto_group_bin_0235 = frame (4k)
frame_crypto_group_bin_0236 = frame (4k)
frame_crypto_group_bin_0237 = frame (4k)
frame_crypto_group_bin_0238 = frame (4k)
frame_crypto_group_bin_0239 = frame (4k)
frame_crypto_group_bin_0240 = frame (4k)
frame_crypto_group_bin_0241 = frame (4k)
frame_crypto_group_bin_0242 = frame (4k)
frame_crypto_group_bin_0243 = frame (4k)
frame_crypto_group_bin_0244 = frame (4k)
frame_crypto_group_bin_0245 = frame (4k)
frame_crypto_group_bin_0246 = frame (4k)
frame_crypto_group_bin_0247 = frame (4k)
frame_crypto_group_bin_0249 = frame (4k)
frame_crypto_group_bin_0250 = frame (4k)
frame_crypto_group_bin_0251 = frame (4k)
frame_crypto_group_bin_0252 = frame (4k)
frame_crypto_group_bin_0253 = frame (4k)
frame_crypto_group_bin_0254 = frame (4k)
frame_crypto_group_bin_0256 = frame (4k)
frame_crypto_group_bin_0257 = frame (4k)
frame_crypto_group_bin_0258 = frame (4k)
frame_crypto_group_bin_0259 = frame (4k)
frame_crypto_group_bin_0260 = frame (4k)
frame_crypto_group_bin_0261 = frame (4k)
frame_crypto_group_bin_0262 = frame (4k)
frame_crypto_group_bin_0263 = frame (4k)
frame_crypto_group_bin_0264 = frame (4k)
frame_crypto_group_bin_0265 = frame (4k)
frame_crypto_group_bin_0266 = frame (4k)
frame_crypto_group_bin_0267 = frame (4k)
frame_crypto_group_bin_0268 = frame (4k)
frame_crypto_group_bin_0269 = frame (4k)
frame_crypto_group_bin_0270 = frame (4k)
frame_crypto_group_bin_0271 = frame (4k)
frame_crypto_group_bin_0272 = frame (4k)
frame_crypto_group_bin_0273 = frame (4k)
frame_crypto_group_bin_0274 = frame (4k)
frame_crypto_group_bin_0275 = frame (4k)
frame_crypto_group_bin_0276 = frame (4k)
frame_crypto_group_bin_0277 = frame (4k)
frame_crypto_group_bin_0278 = frame (4k)
frame_crypto_group_bin_0279 = frame (4k)
frame_crypto_group_bin_0280 = frame (4k)
frame_crypto_group_bin_0281 = frame (4k)
frame_crypto_group_bin_0282 = frame (4k)
frame_crypto_group_bin_0283 = frame (4k)
frame_crypto_group_bin_0284 = frame (4k)
frame_crypto_group_bin_0285 = frame (4k)
frame_crypto_group_bin_0286 = frame (4k)
frame_crypto_group_bin_0287 = frame (4k)
frame_crypto_group_bin_0289 = frame (4k)
frame_crypto_group_bin_0290 = frame (4k)
frame_crypto_group_bin_0291 = frame (4k)
frame_crypto_group_bin_0292 = frame (4k)
frame_crypto_group_bin_0293 = frame (4k)
frame_crypto_group_bin_0294 = frame (4k)
frame_crypto_group_bin_0295 = frame (4k)
frame_crypto_group_bin_0296 = frame (4k)
frame_crypto_group_bin_0297 = frame (4k)
frame_crypto_group_bin_0298 = frame (4k)
frame_crypto_group_bin_0299 = frame (4k)
frame_crypto_group_bin_0300 = frame (4k)
frame_crypto_group_bin_0301 = frame (4k)
frame_crypto_group_bin_0302 = frame (4k)
frame_crypto_group_bin_0304 = frame (4k)
frame_crypto_group_bin_0305 = frame (4k)
frame_crypto_group_bin_0306 = frame (4k)
frame_crypto_group_bin_0307 = frame (4k)
frame_crypto_group_bin_0308 = frame (4k)
frame_crypto_group_bin_0309 = frame (4k)
frame_crypto_group_bin_0310 = frame (4k)
frame_crypto_group_bin_0311 = frame (4k)
frame_crypto_group_bin_0312 = frame (4k)
frame_crypto_group_bin_0313 = frame (4k)
frame_crypto_group_bin_0314 = frame (4k)
frame_crypto_group_bin_0315 = frame (4k)
frame_crypto_group_bin_0317 = frame (4k)
frame_crypto_group_bin_0319 = frame (4k)
frame_crypto_group_bin_0320 = frame (4k)
frame_crypto_group_bin_0321 = frame (4k)
frame_crypto_group_bin_0322 = frame (4k)
frame_crypto_group_bin_0323 = frame (4k)
frame_crypto_group_bin_0324 = frame (4k)
frame_modchk_group_bin_0000 = frame (4k)
frame_modchk_group_bin_0001 = frame (4k)
frame_modchk_group_bin_0002 = frame (4k)
frame_modchk_group_bin_0003 = frame (4k)
frame_modchk_group_bin_0004 = frame (4k)
frame_modchk_group_bin_0005 = frame (4k)
frame_modchk_group_bin_0006 = frame (4k)
frame_modchk_group_bin_0007 = frame (4k)
frame_modchk_group_bin_0008 = frame (4k)
frame_modchk_group_bin_0010 = frame (4k)
frame_modchk_group_bin_0011 = frame (4k)
frame_modchk_group_bin_0012 = frame (4k)
frame_modchk_group_bin_0013 = frame (4k)
frame_modchk_group_bin_0014 = frame (4k)
frame_modchk_group_bin_0015 = frame (4k)
frame_modchk_group_bin_0016 = frame (4k)
frame_modchk_group_bin_0017 = frame (4k)
frame_modchk_group_bin_0018 = frame (4k)
frame_modchk_group_bin_0019 = frame (4k)
frame_modchk_group_bin_0020 = frame (4k)
frame_modchk_group_bin_0021 = frame (4k)
frame_modchk_group_bin_0022 = frame (4k)
frame_modchk_group_bin_0023 = frame (4k)
frame_modchk_group_bin_0024 = frame (4k)
frame_modchk_group_bin_0025 = frame (4k)
frame_modchk_group_bin_0026 = frame (4k)
frame_modchk_group_bin_0027 = frame (4k)
frame_modchk_group_bin_0028 = frame (4k)
frame_modchk_group_bin_0029 = frame (4k)
frame_modchk_group_bin_0030 = frame (4k)
frame_modchk_group_bin_0031 = frame (4k)
frame_modchk_group_bin_0032 = frame (4k)
frame_modchk_group_bin_0035 = frame (4k)
frame_modchk_group_bin_0037 = frame (4k)
frame_modchk_group_bin_0038 = frame (4k)
frame_modchk_group_bin_0039 = frame (4k)
frame_modchk_group_bin_0041 = frame (4k)
frame_modchk_group_bin_0042 = frame (4k)
frame_modchk_group_bin_0043 = frame (4k)
frame_modchk_group_bin_0044 = frame (4k)
frame_modchk_group_bin_0045 = frame (4k)
frame_modchk_group_bin_0046 = frame (4k)
frame_modchk_group_bin_0047 = frame (4k)
frame_modchk_group_bin_0048 = frame (4k)
frame_modchk_group_bin_0049 = frame (4k)
frame_modchk_group_bin_0051 = frame (4k)
frame_modchk_group_bin_0052 = frame (4k)
frame_modchk_group_bin_0053 = frame (4k)
frame_modchk_group_bin_0054 = frame (4k)
frame_modchk_group_bin_0055 = frame (4k)
frame_modchk_group_bin_0056 = frame (4k)
frame_modchk_group_bin_0057 = frame (4k)
frame_modchk_group_bin_0058 = frame (4k)
frame_modchk_group_bin_0059 = frame (4k)
frame_modchk_group_bin_0060 = frame (4k)
frame_modchk_group_bin_0061 = frame (4k)
frame_modchk_group_bin_0062 = frame (4k)
frame_modchk_group_bin_0063 = frame (4k)
frame_modchk_group_bin_0065 = frame (4k)
frame_modchk_group_bin_0067 = frame (4k)
frame_modchk_group_bin_0068 = frame (4k)
frame_modchk_group_bin_0070 = frame (4k)
frame_modchk_group_bin_0071 = frame (4k)
frame_modchk_group_bin_0072 = frame (4k)
frame_modchk_group_bin_0073 = frame (4k)
frame_modchk_group_bin_0074 = frame (4k)
frame_modchk_group_bin_0075 = frame (4k)
frame_modchk_group_bin_0076 = frame (4k)
frame_modchk_group_bin_0077 = frame (4k)
frame_modchk_group_bin_0078 = frame (4k)
frame_modchk_group_bin_0080 = frame (4k)
frame_modchk_group_bin_0081 = frame (4k)
frame_modchk_group_bin_0083 = frame (4k)
frame_modchk_group_bin_0084 = frame (4k)
frame_modchk_group_bin_0085 = frame (4k)
frame_modchk_group_bin_0086 = frame (4k)
frame_modchk_group_bin_0087 = frame (4k)
frame_modchk_group_bin_0088 = frame (4k)
frame_modchk_group_bin_0089 = frame (4k)
frame_modchk_group_bin_0090 = frame (4k)
frame_modchk_group_bin_0091 = frame (4k)
frame_modchk_group_bin_0092 = frame (4k)
frame_modchk_group_bin_0093 = frame (4k)
frame_modchk_group_bin_0094 = frame (4k)
frame_modchk_group_bin_0095 = frame (4k)
frame_modchk_group_bin_0096 = frame (4k)
frame_modchk_group_bin_0097 = frame (4k)
frame_modchk_group_bin_0098 = frame (4k)
frame_modchk_group_bin_0099 = frame (4k)
frame_modchk_group_bin_0100 = frame (4k)
frame_modchk_group_bin_0101 = frame (4k)
frame_modchk_group_bin_0102 = frame (4k)
frame_modchk_group_bin_0104 = frame (4k)
frame_modchk_group_bin_0105 = frame (4k)
frame_modchk_group_bin_0106 = frame (4k)
frame_modchk_group_bin_0107 = frame (4k)
frame_modchk_group_bin_0108 = frame (4k)
frame_modchk_group_bin_0109 = frame (4k)
frame_modchk_group_bin_0111 = frame (4k)
frame_modchk_group_bin_0112 = frame (4k)
frame_modchk_group_bin_0114 = frame (4k)
frame_modchk_group_bin_0115 = frame (4k)
frame_modchk_group_bin_0116 = frame (4k)
frame_modchk_group_bin_0117 = frame (4k)
frame_modchk_group_bin_0118 = frame (4k)
frame_modchk_group_bin_0119 = frame (4k)
frame_modchk_group_bin_0120 = frame (4k)
frame_modchk_group_bin_0121 = frame (4k)
frame_modchk_group_bin_0122 = frame (4k)
frame_modchk_group_bin_0123 = frame (4k)
frame_modchk_group_bin_0124 = frame (4k)
frame_modchk_group_bin_0125 = frame (4k)
frame_modchk_group_bin_0126 = frame (4k)
frame_modchk_group_bin_0127 = frame (4k)
frame_modchk_group_bin_0128 = frame (4k)
frame_modchk_group_bin_0129 = frame (4k)
frame_modchk_group_bin_0130 = frame (4k)
frame_modchk_group_bin_0131 = frame (4k)
frame_modchk_group_bin_0132 = frame (4k)
frame_modchk_group_bin_0133 = frame (4k)
frame_modchk_group_bin_0134 = frame (4k)
frame_modchk_group_bin_0136 = frame (4k)
frame_modchk_group_bin_0137 = frame (4k)
frame_modchk_group_bin_0138 = frame (4k)
frame_modchk_group_bin_0139 = frame (4k)
frame_modchk_group_bin_0140 = frame (4k)
frame_modchk_group_bin_0141 = frame (4k)
frame_modchk_group_bin_0142 = frame (4k)
frame_modchk_group_bin_0143 = frame (4k)
frame_modchk_group_bin_0144 = frame (4k)
frame_modchk_group_bin_0145 = frame (4k)
frame_modchk_group_bin_0146 = frame (4k)
frame_modchk_group_bin_0147 = frame (4k)
frame_modchk_group_bin_0148 = frame (4k)
frame_modchk_group_bin_0149 = frame (4k)
frame_modchk_group_bin_0150 = frame (4k)
frame_modchk_group_bin_0151 = frame (4k)
frame_modchk_group_bin_0152 = frame (4k)
frame_modchk_group_bin_0153 = frame (4k)
frame_modchk_group_bin_0154 = frame (4k)
frame_modchk_group_bin_0155 = frame (4k)
frame_modchk_group_bin_0157 = frame (4k)
frame_modchk_group_bin_0158 = frame (4k)
frame_modchk_group_bin_0159 = frame (4k)
frame_modchk_group_bin_0160 = frame (4k)
frame_modchk_group_bin_0161 = frame (4k)
frame_modchk_group_bin_0162 = frame (4k)
frame_modchk_group_bin_0163 = frame (4k)
frame_modchk_group_bin_0164 = frame (4k)
frame_modchk_group_bin_0165 = frame (4k)
frame_modchk_group_bin_0166 = frame (4k)
frame_modchk_group_bin_0167 = frame (4k)
frame_modchk_group_bin_0168 = frame (4k)
frame_modchk_group_bin_0169 = frame (4k)
frame_modchk_group_bin_0170 = frame (4k)
frame_modchk_group_bin_0171 = frame (4k)
frame_modchk_group_bin_0173 = frame (4k)
frame_modchk_group_bin_0174 = frame (4k)
frame_modchk_group_bin_0176 = frame (4k)
frame_modchk_group_bin_0177 = frame (4k)
frame_modchk_group_bin_0178 = frame (4k)
frame_modchk_group_bin_0179 = frame (4k)
frame_modchk_group_bin_0180 = frame (4k)
frame_modchk_group_bin_0181 = frame (4k)
frame_modchk_group_bin_0183 = frame (4k)
frame_modchk_group_bin_0184 = frame (4k)
frame_modchk_group_bin_0185 = frame (4k)
frame_modchk_group_bin_0186 = frame (4k)
frame_modchk_group_bin_0187 = frame (4k)
frame_modchk_group_bin_0188 = frame (4k)
frame_modchk_group_bin_0189 = frame (4k)
frame_modchk_group_bin_0190 = frame (4k)
frame_modchk_group_bin_0191 = frame (4k)
frame_modchk_group_bin_0192 = frame (4k)
frame_modchk_group_bin_0193 = frame (4k)
frame_modchk_group_bin_0194 = frame (4k)
frame_modchk_group_bin_0195 = frame (4k)
frame_modchk_group_bin_0196 = frame (4k)
frame_modchk_group_bin_0197 = frame (4k)
frame_modchk_group_bin_0198 = frame (4k)
frame_modchk_group_bin_0199 = frame (4k)
frame_modchk_group_bin_0200 = frame (4k)
frame_modchk_group_bin_0201 = frame (4k)
frame_modchk_group_bin_0202 = frame (4k)
frame_modchk_group_bin_0203 = frame (4k)
frame_modchk_group_bin_0204 = frame (4k)
frame_modchk_group_bin_0205 = frame (4k)
frame_modchk_group_bin_0206 = frame (4k)
frame_modchk_group_bin_0207 = frame (4k)
frame_modchk_group_bin_0208 = frame (4k)
frame_modchk_group_bin_0209 = frame (4k)
frame_modchk_group_bin_0210 = frame (4k)
frame_modchk_group_bin_0211 = frame (4k)
frame_modchk_group_bin_0212 = frame (4k)
frame_modchk_group_bin_0213 = frame (4k)
frame_modchk_group_bin_0214 = frame (4k)
frame_modchk_group_bin_0215 = frame (4k)
frame_modchk_group_bin_0216 = frame (4k)
frame_modchk_group_bin_0217 = frame (4k)
frame_modchk_group_bin_0218 = frame (4k)
frame_modchk_group_bin_0220 = frame (4k)
frame_modchk_group_bin_0221 = frame (4k)
frame_modchk_group_bin_0222 = frame (4k)
frame_modchk_group_bin_0223 = frame (4k)
frame_modchk_group_bin_0224 = frame (4k)
frame_modchk_group_bin_0225 = frame (4k)
frame_modchk_group_bin_0226 = frame (4k)
frame_modchk_group_bin_0228 = frame (4k)
frame_modchk_group_bin_0229 = frame (4k)
frame_modchk_group_bin_0230 = frame (4k)
frame_modchk_group_bin_0231 = frame (4k)
frame_modchk_group_bin_0232 = frame (4k)
frame_modchk_group_bin_0233 = frame (4k)
frame_modchk_group_bin_0234 = frame (4k)
frame_modchk_group_bin_0235 = frame (4k)
frame_modchk_group_bin_0236 = frame (4k)
frame_modchk_group_bin_0237 = frame (4k)
frame_modchk_group_bin_0238 = frame (4k)
frame_modchk_group_bin_0239 = frame (4k)
frame_modchk_group_bin_0240 = frame (4k)
frame_modchk_group_bin_0241 = frame (4k)
frame_modchk_group_bin_0242 = frame (4k)
frame_modchk_group_bin_0243 = frame (4k)
frame_modchk_group_bin_0244 = frame (4k)
frame_modchk_group_bin_0245 = frame (4k)
frame_modchk_group_bin_0246 = frame (4k)
frame_modchk_group_bin_0248 = frame (4k)
frame_modchk_group_bin_0249 = frame (4k)
frame_modchk_group_bin_0250 = frame (4k)
frame_modchk_group_bin_0251 = frame (4k)
frame_modchk_group_bin_0252 = frame (4k)
frame_modchk_group_bin_0253 = frame (4k)
frame_modchk_group_bin_0255 = frame (4k)
frame_modchk_group_bin_0256 = frame (4k)
frame_modchk_group_bin_0257 = frame (4k)
frame_modchk_group_bin_0258 = frame (4k)
frame_modchk_group_bin_0259 = frame (4k)
frame_modchk_group_bin_0260 = frame (4k)
frame_modchk_group_bin_0261 = frame (4k)
frame_modchk_group_bin_0262 = frame (4k)
frame_modchk_group_bin_0263 = frame (4k)
frame_modchk_group_bin_0264 = frame (4k)
frame_modchk_group_bin_0265 = frame (4k)
frame_modchk_group_bin_0266 = frame (4k)
frame_modchk_group_bin_0267 = frame (4k)
frame_modchk_group_bin_0268 = frame (4k)
frame_modchk_group_bin_0269 = frame (4k)
frame_modchk_group_bin_0270 = frame (4k)
frame_modchk_group_bin_0271 = frame (4k)
frame_modchk_group_bin_0272 = frame (4k)
frame_modchk_group_bin_0273 = frame (4k)
frame_modchk_group_bin_0274 = frame (4k)
frame_modchk_group_bin_0275 = frame (4k)
frame_modchk_group_bin_0276 = frame (4k)
frame_modchk_group_bin_0277 = frame (4k)
frame_modchk_group_bin_0278 = frame (4k)
frame_modchk_group_bin_0279 = frame (4k)
frame_modchk_group_bin_0280 = frame (4k)
frame_modchk_group_bin_0281 = frame (4k)
frame_modchk_group_bin_0282 = frame (4k)
frame_modchk_group_bin_0283 = frame (4k)
frame_modchk_group_bin_0284 = frame (4k)
frame_modchk_group_bin_0285 = frame (4k)
frame_modchk_group_bin_0286 = frame (4k)
frame_modchk_group_bin_0288 = frame (4k)
frame_modchk_group_bin_0289 = frame (4k)
frame_modchk_group_bin_0290 = frame (4k)
frame_modchk_group_bin_0291 = frame (4k)
frame_modchk_group_bin_0292 = frame (4k)
frame_modchk_group_bin_0293 = frame (4k)
frame_modchk_group_bin_0294 = frame (4k)
frame_modchk_group_bin_0295 = frame (4k)
frame_modchk_group_bin_0296 = frame (4k)
frame_modchk_group_bin_0297 = frame (4k)
frame_modchk_group_bin_0298 = frame (4k)
frame_modchk_group_bin_0299 = frame (4k)
frame_modchk_group_bin_0300 = frame (4k)
frame_modchk_group_bin_0301 = frame (4k)
frame_modchk_group_bin_0303 = frame (4k)
frame_modchk_group_bin_0304 = frame (4k)
frame_modchk_group_bin_0305 = frame (4k)
frame_modchk_group_bin_0306 = frame (4k)
frame_modchk_group_bin_0307 = frame (4k)
frame_modchk_group_bin_0308 = frame (4k)
frame_modchk_group_bin_0309 = frame (4k)
frame_modchk_group_bin_0310 = frame (4k)
frame_modchk_group_bin_0311 = frame (4k)
frame_modchk_group_bin_0312 = frame (4k)
frame_modchk_group_bin_0313 = frame (4k)
frame_modchk_group_bin_0314 = frame (4k)
frame_modchk_group_bin_0316 = frame (4k)
frame_modchk_group_bin_0318 = frame (4k)
frame_modchk_group_bin_0319 = frame (4k)
frame_modchk_group_bin_0320 = frame (4k)
frame_modchk_group_bin_0321 = frame (4k)
frame_modchk_group_bin_0322 = frame (4k)
frame_modchk_group_bin_0323 = frame (4k)
frame_modtx_group_bin_0000 = frame (4k)
frame_modtx_group_bin_0001 = frame (4k)
frame_modtx_group_bin_0002 = frame (4k)
frame_modtx_group_bin_0003 = frame (4k)
frame_modtx_group_bin_0004 = frame (4k)
frame_modtx_group_bin_0005 = frame (4k)
frame_modtx_group_bin_0006 = frame (4k)
frame_modtx_group_bin_0007 = frame (4k)
frame_modtx_group_bin_0008 = frame (4k)
frame_modtx_group_bin_0010 = frame (4k)
frame_modtx_group_bin_0011 = frame (4k)
frame_modtx_group_bin_0012 = frame (4k)
frame_modtx_group_bin_0013 = frame (4k)
frame_modtx_group_bin_0014 = frame (4k)
frame_modtx_group_bin_0015 = frame (4k)
frame_modtx_group_bin_0016 = frame (4k)
frame_modtx_group_bin_0017 = frame (4k)
frame_modtx_group_bin_0018 = frame (4k)
frame_modtx_group_bin_0019 = frame (4k)
frame_modtx_group_bin_0020 = frame (4k)
frame_modtx_group_bin_0021 = frame (4k)
frame_modtx_group_bin_0022 = frame (4k)
frame_modtx_group_bin_0023 = frame (4k)
frame_modtx_group_bin_0024 = frame (4k)
frame_modtx_group_bin_0025 = frame (4k)
frame_modtx_group_bin_0026 = frame (4k)
frame_modtx_group_bin_0027 = frame (4k)
frame_modtx_group_bin_0028 = frame (4k)
frame_modtx_group_bin_0029 = frame (4k)
frame_modtx_group_bin_0030 = frame (4k)
frame_modtx_group_bin_0031 = frame (4k)
frame_modtx_group_bin_0032 = frame (4k)
frame_modtx_group_bin_0035 = frame (4k)
frame_modtx_group_bin_0037 = frame (4k)
frame_modtx_group_bin_0038 = frame (4k)
frame_modtx_group_bin_0039 = frame (4k)
frame_modtx_group_bin_0041 = frame (4k)
frame_modtx_group_bin_0042 = frame (4k)
frame_modtx_group_bin_0043 = frame (4k)
frame_modtx_group_bin_0044 = frame (4k)
frame_modtx_group_bin_0045 = frame (4k)
frame_modtx_group_bin_0046 = frame (4k)
frame_modtx_group_bin_0047 = frame (4k)
frame_modtx_group_bin_0048 = frame (4k)
frame_modtx_group_bin_0049 = frame (4k)
frame_modtx_group_bin_0051 = frame (4k)
frame_modtx_group_bin_0052 = frame (4k)
frame_modtx_group_bin_0053 = frame (4k)
frame_modtx_group_bin_0054 = frame (4k)
frame_modtx_group_bin_0055 = frame (4k)
frame_modtx_group_bin_0056 = frame (4k)
frame_modtx_group_bin_0057 = frame (4k)
frame_modtx_group_bin_0058 = frame (4k)
frame_modtx_group_bin_0059 = frame (4k)
frame_modtx_group_bin_0060 = frame (4k)
frame_modtx_group_bin_0061 = frame (4k)
frame_modtx_group_bin_0062 = frame (4k)
frame_modtx_group_bin_0063 = frame (4k)
frame_modtx_group_bin_0065 = frame (4k)
frame_modtx_group_bin_0067 = frame (4k)
frame_modtx_group_bin_0068 = frame (4k)
frame_modtx_group_bin_0070 = frame (4k)
frame_modtx_group_bin_0071 = frame (4k)
frame_modtx_group_bin_0072 = frame (4k)
frame_modtx_group_bin_0073 = frame (4k)
frame_modtx_group_bin_0074 = frame (4k)
frame_modtx_group_bin_0075 = frame (4k)
frame_modtx_group_bin_0076 = frame (4k)
frame_modtx_group_bin_0077 = frame (4k)
frame_modtx_group_bin_0078 = frame (4k)
frame_modtx_group_bin_0080 = frame (4k)
frame_modtx_group_bin_0081 = frame (4k)
frame_modtx_group_bin_0083 = frame (4k)
frame_modtx_group_bin_0084 = frame (4k)
frame_modtx_group_bin_0085 = frame (4k)
frame_modtx_group_bin_0086 = frame (4k)
frame_modtx_group_bin_0087 = frame (4k)
frame_modtx_group_bin_0088 = frame (4k)
frame_modtx_group_bin_0089 = frame (4k)
frame_modtx_group_bin_0090 = frame (4k)
frame_modtx_group_bin_0091 = frame (4k)
frame_modtx_group_bin_0092 = frame (4k)
frame_modtx_group_bin_0093 = frame (4k)
frame_modtx_group_bin_0094 = frame (4k)
frame_modtx_group_bin_0095 = frame (4k)
frame_modtx_group_bin_0096 = frame (4k)
frame_modtx_group_bin_0097 = frame (4k)
frame_modtx_group_bin_0098 = frame (4k)
frame_modtx_group_bin_0099 = frame (4k)
frame_modtx_group_bin_0100 = frame (4k)
frame_modtx_group_bin_0101 = frame (4k)
frame_modtx_group_bin_0102 = frame (4k)
frame_modtx_group_bin_0104 = frame (4k)
frame_modtx_group_bin_0105 = frame (4k)
frame_modtx_group_bin_0106 = frame (4k)
frame_modtx_group_bin_0107 = frame (4k)
frame_modtx_group_bin_0108 = frame (4k)
frame_modtx_group_bin_0109 = frame (4k)
frame_modtx_group_bin_0111 = frame (4k)
frame_modtx_group_bin_0112 = frame (4k)
frame_modtx_group_bin_0114 = frame (4k)
frame_modtx_group_bin_0115 = frame (4k)
frame_modtx_group_bin_0116 = frame (4k)
frame_modtx_group_bin_0117 = frame (4k)
frame_modtx_group_bin_0118 = frame (4k)
frame_modtx_group_bin_0119 = frame (4k)
frame_modtx_group_bin_0120 = frame (4k)
frame_modtx_group_bin_0121 = frame (4k)
frame_modtx_group_bin_0122 = frame (4k)
frame_modtx_group_bin_0123 = frame (4k)
frame_modtx_group_bin_0124 = frame (4k)
frame_modtx_group_bin_0125 = frame (4k)
frame_modtx_group_bin_0126 = frame (4k)
frame_modtx_group_bin_0127 = frame (4k)
frame_modtx_group_bin_0128 = frame (4k)
frame_modtx_group_bin_0129 = frame (4k)
frame_modtx_group_bin_0130 = frame (4k)
frame_modtx_group_bin_0131 = frame (4k)
frame_modtx_group_bin_0132 = frame (4k)
frame_modtx_group_bin_0133 = frame (4k)
frame_modtx_group_bin_0134 = frame (4k)
frame_modtx_group_bin_0136 = frame (4k)
frame_modtx_group_bin_0137 = frame (4k)
frame_modtx_group_bin_0138 = frame (4k)
frame_modtx_group_bin_0139 = frame (4k)
frame_modtx_group_bin_0140 = frame (4k)
frame_modtx_group_bin_0141 = frame (4k)
frame_modtx_group_bin_0142 = frame (4k)
frame_modtx_group_bin_0143 = frame (4k)
frame_modtx_group_bin_0144 = frame (4k)
frame_modtx_group_bin_0145 = frame (4k)
frame_modtx_group_bin_0146 = frame (4k)
frame_modtx_group_bin_0147 = frame (4k)
frame_modtx_group_bin_0148 = frame (4k)
frame_modtx_group_bin_0149 = frame (4k)
frame_modtx_group_bin_0150 = frame (4k)
frame_modtx_group_bin_0151 = frame (4k)
frame_modtx_group_bin_0152 = frame (4k)
frame_modtx_group_bin_0153 = frame (4k)
frame_modtx_group_bin_0154 = frame (4k)
frame_modtx_group_bin_0155 = frame (4k)
frame_modtx_group_bin_0157 = frame (4k)
frame_modtx_group_bin_0158 = frame (4k)
frame_modtx_group_bin_0159 = frame (4k)
frame_modtx_group_bin_0160 = frame (4k)
frame_modtx_group_bin_0161 = frame (4k)
frame_modtx_group_bin_0162 = frame (4k)
frame_modtx_group_bin_0163 = frame (4k)
frame_modtx_group_bin_0164 = frame (4k)
frame_modtx_group_bin_0165 = frame (4k)
frame_modtx_group_bin_0166 = frame (4k)
frame_modtx_group_bin_0167 = frame (4k)
frame_modtx_group_bin_0168 = frame (4k)
frame_modtx_group_bin_0169 = frame (4k)
frame_modtx_group_bin_0170 = frame (4k)
frame_modtx_group_bin_0171 = frame (4k)
frame_modtx_group_bin_0172 = frame (4k)
frame_modtx_group_bin_0173 = frame (4k)
frame_modtx_group_bin_0175 = frame (4k)
frame_modtx_group_bin_0176 = frame (4k)
frame_modtx_group_bin_0177 = frame (4k)
frame_modtx_group_bin_0178 = frame (4k)
frame_modtx_group_bin_0179 = frame (4k)
frame_modtx_group_bin_0180 = frame (4k)
frame_modtx_group_bin_0182 = frame (4k)
frame_modtx_group_bin_0183 = frame (4k)
frame_modtx_group_bin_0184 = frame (4k)
frame_modtx_group_bin_0185 = frame (4k)
frame_modtx_group_bin_0186 = frame (4k)
frame_modtx_group_bin_0187 = frame (4k)
frame_modtx_group_bin_0188 = frame (4k)
frame_modtx_group_bin_0189 = frame (4k)
frame_modtx_group_bin_0190 = frame (4k)
frame_modtx_group_bin_0191 = frame (4k)
frame_modtx_group_bin_0192 = frame (4k)
frame_modtx_group_bin_0193 = frame (4k)
frame_modtx_group_bin_0194 = frame (4k)
frame_modtx_group_bin_0195 = frame (4k)
frame_modtx_group_bin_0196 = frame (4k)
frame_modtx_group_bin_0197 = frame (4k)
frame_modtx_group_bin_0198 = frame (4k)
frame_modtx_group_bin_0199 = frame (4k)
frame_modtx_group_bin_0200 = frame (4k)
frame_modtx_group_bin_0201 = frame (4k)
frame_modtx_group_bin_0202 = frame (4k)
frame_modtx_group_bin_0203 = frame (4k)
frame_modtx_group_bin_0204 = frame (4k)
frame_modtx_group_bin_0205 = frame (4k)
frame_modtx_group_bin_0206 = frame (4k)
frame_modtx_group_bin_0207 = frame (4k)
frame_modtx_group_bin_0208 = frame (4k)
frame_modtx_group_bin_0209 = frame (4k)
frame_modtx_group_bin_0210 = frame (4k)
frame_modtx_group_bin_0211 = frame (4k)
frame_modtx_group_bin_0212 = frame (4k)
frame_modtx_group_bin_0213 = frame (4k)
frame_modtx_group_bin_0214 = frame (4k)
frame_modtx_group_bin_0215 = frame (4k)
frame_modtx_group_bin_0216 = frame (4k)
frame_modtx_group_bin_0217 = frame (4k)
frame_modtx_group_bin_0219 = frame (4k)
frame_modtx_group_bin_0220 = frame (4k)
frame_modtx_group_bin_0221 = frame (4k)
frame_modtx_group_bin_0222 = frame (4k)
frame_modtx_group_bin_0223 = frame (4k)
frame_modtx_group_bin_0224 = frame (4k)
frame_modtx_group_bin_0225 = frame (4k)
frame_modtx_group_bin_0227 = frame (4k)
frame_modtx_group_bin_0228 = frame (4k)
frame_modtx_group_bin_0229 = frame (4k)
frame_modtx_group_bin_0230 = frame (4k)
frame_modtx_group_bin_0231 = frame (4k)
frame_modtx_group_bin_0232 = frame (4k)
frame_modtx_group_bin_0233 = frame (4k)
frame_modtx_group_bin_0234 = frame (4k)
frame_modtx_group_bin_0235 = frame (4k)
frame_modtx_group_bin_0236 = frame (4k)
frame_modtx_group_bin_0237 = frame (4k)
frame_modtx_group_bin_0238 = frame (4k)
frame_modtx_group_bin_0239 = frame (4k)
frame_modtx_group_bin_0240 = frame (4k)
frame_modtx_group_bin_0241 = frame (4k)
frame_modtx_group_bin_0242 = frame (4k)
frame_modtx_group_bin_0243 = frame (4k)
frame_modtx_group_bin_0244 = frame (4k)
frame_modtx_group_bin_0245 = frame (4k)
frame_modtx_group_bin_0247 = frame (4k)
frame_modtx_group_bin_0248 = frame (4k)
frame_modtx_group_bin_0249 = frame (4k)
frame_modtx_group_bin_0250 = frame (4k)
frame_modtx_group_bin_0251 = frame (4k)
frame_modtx_group_bin_0252 = frame (4k)
frame_modtx_group_bin_0254 = frame (4k)
frame_modtx_group_bin_0255 = frame (4k)
frame_modtx_group_bin_0256 = frame (4k)
frame_modtx_group_bin_0257 = frame (4k)
frame_modtx_group_bin_0259 = frame (4k)
frame_modtx_group_bin_0260 = frame (4k)
frame_modtx_group_bin_0261 = frame (4k)
frame_modtx_group_bin_0262 = frame (4k)
frame_modtx_group_bin_0263 = frame (4k)
frame_modtx_group_bin_0264 = frame (4k)
frame_modtx_group_bin_0265 = frame (4k)
frame_modtx_group_bin_0266 = frame (4k)
frame_modtx_group_bin_0267 = frame (4k)
frame_modtx_group_bin_0268 = frame (4k)
frame_modtx_group_bin_0269 = frame (4k)
frame_modtx_group_bin_0270 = frame (4k)
frame_modtx_group_bin_0271 = frame (4k)
frame_modtx_group_bin_0272 = frame (4k)
frame_modtx_group_bin_0273 = frame (4k)
frame_modtx_group_bin_0274 = frame (4k)
frame_modtx_group_bin_0275 = frame (4k)
frame_modtx_group_bin_0276 = frame (4k)
frame_modtx_group_bin_0277 = frame (4k)
frame_modtx_group_bin_0278 = frame (4k)
frame_modtx_group_bin_0279 = frame (4k)
frame_modtx_group_bin_0280 = frame (4k)
frame_modtx_group_bin_0281 = frame (4k)
frame_modtx_group_bin_0282 = frame (4k)
frame_modtx_group_bin_0283 = frame (4k)
frame_modtx_group_bin_0284 = frame (4k)
frame_modtx_group_bin_0285 = frame (4k)
frame_modtx_group_bin_0287 = frame (4k)
frame_modtx_group_bin_0288 = frame (4k)
frame_modtx_group_bin_0289 = frame (4k)
frame_modtx_group_bin_0290 = frame (4k)
frame_modtx_group_bin_0291 = frame (4k)
frame_modtx_group_bin_0292 = frame (4k)
frame_modtx_group_bin_0293 = frame (4k)
frame_modtx_group_bin_0294 = frame (4k)
frame_modtx_group_bin_0295 = frame (4k)
frame_modtx_group_bin_0296 = frame (4k)
frame_modtx_group_bin_0297 = frame (4k)
frame_modtx_group_bin_0298 = frame (4k)
frame_modtx_group_bin_0299 = frame (4k)
frame_modtx_group_bin_0300 = frame (4k)
frame_modtx_group_bin_0302 = frame (4k)
frame_modtx_group_bin_0303 = frame (4k)
frame_modtx_group_bin_0304 = frame (4k)
frame_modtx_group_bin_0305 = frame (4k)
frame_modtx_group_bin_0306 = frame (4k)
frame_modtx_group_bin_0307 = frame (4k)
frame_modtx_group_bin_0308 = frame (4k)
frame_modtx_group_bin_0309 = frame (4k)
frame_modtx_group_bin_0310 = frame (4k)
frame_modtx_group_bin_0311 = frame (4k)
frame_modtx_group_bin_0312 = frame (4k)
frame_modtx_group_bin_0313 = frame (4k)
frame_modtx_group_bin_0315 = frame (4k)
frame_modtx_group_bin_0317 = frame (4k)
frame_modtx_group_bin_0318 = frame (4k)
frame_modtx_group_bin_0319 = frame (4k)
frame_modtx_group_bin_0320 = frame (4k)
frame_modtx_group_bin_0321 = frame (4k)
frame_modtx_group_bin_0322 = frame (4k)
frame_signtx_group_bin_0000 = frame (4k)
frame_signtx_group_bin_0001 = frame (4k)
frame_signtx_group_bin_0002 = frame (4k)
frame_signtx_group_bin_0003 = frame (4k)
frame_signtx_group_bin_0004 = frame (4k)
frame_signtx_group_bin_0005 = frame (4k)
frame_signtx_group_bin_0006 = frame (4k)
frame_signtx_group_bin_0007 = frame (4k)
frame_signtx_group_bin_0008 = frame (4k)
frame_signtx_group_bin_0009 = frame (4k)
frame_signtx_group_bin_0010 = frame (4k)
frame_signtx_group_bin_0011 = frame (4k)
frame_signtx_group_bin_0012 = frame (4k)
frame_signtx_group_bin_0013 = frame (4k)
frame_signtx_group_bin_0014 = frame (4k)
frame_signtx_group_bin_0015 = frame (4k)
frame_signtx_group_bin_0016 = frame (4k)
frame_signtx_group_bin_0017 = frame (4k)
frame_signtx_group_bin_0018 = frame (4k)
frame_signtx_group_bin_0019 = frame (4k)
frame_signtx_group_bin_0020 = frame (4k)
frame_signtx_group_bin_0021 = frame (4k)
frame_signtx_group_bin_0022 = frame (4k)
frame_signtx_group_bin_0023 = frame (4k)
frame_signtx_group_bin_0024 = frame (4k)
frame_signtx_group_bin_0025 = frame (4k)
frame_signtx_group_bin_0026 = frame (4k)
frame_signtx_group_bin_0027 = frame (4k)
frame_signtx_group_bin_0028 = frame (4k)
frame_signtx_group_bin_0029 = frame (4k)
frame_signtx_group_bin_0030 = frame (4k)
frame_signtx_group_bin_0031 = frame (4k)
frame_signtx_group_bin_0032 = frame (4k)
frame_signtx_group_bin_0035 = frame (4k)
frame_signtx_group_bin_0037 = frame (4k)
frame_signtx_group_bin_0038 = frame (4k)
frame_signtx_group_bin_0039 = frame (4k)
frame_signtx_group_bin_0041 = frame (4k)
frame_signtx_group_bin_0042 = frame (4k)
frame_signtx_group_bin_0043 = frame (4k)
frame_signtx_group_bin_0044 = frame (4k)
frame_signtx_group_bin_0045 = frame (4k)
frame_signtx_group_bin_0046 = frame (4k)
frame_signtx_group_bin_0047 = frame (4k)
frame_signtx_group_bin_0048 = frame (4k)
frame_signtx_group_bin_0049 = frame (4k)
frame_signtx_group_bin_0051 = frame (4k)
frame_signtx_group_bin_0052 = frame (4k)
frame_signtx_group_bin_0053 = frame (4k)
frame_signtx_group_bin_0054 = frame (4k)
frame_signtx_group_bin_0055 = frame (4k)
frame_signtx_group_bin_0056 = frame (4k)
frame_signtx_group_bin_0057 = frame (4k)
frame_signtx_group_bin_0058 = frame (4k)
frame_signtx_group_bin_0059 = frame (4k)
frame_signtx_group_bin_0060 = frame (4k)
frame_signtx_group_bin_0061 = frame (4k)
frame_signtx_group_bin_0062 = frame (4k)
frame_signtx_group_bin_0063 = frame (4k)
frame_signtx_group_bin_0065 = frame (4k)
frame_signtx_group_bin_0067 = frame (4k)
frame_signtx_group_bin_0068 = frame (4k)
frame_signtx_group_bin_0070 = frame (4k)
frame_signtx_group_bin_0071 = frame (4k)
frame_signtx_group_bin_0072 = frame (4k)
frame_signtx_group_bin_0073 = frame (4k)
frame_signtx_group_bin_0074 = frame (4k)
frame_signtx_group_bin_0075 = frame (4k)
frame_signtx_group_bin_0076 = frame (4k)
frame_signtx_group_bin_0077 = frame (4k)
frame_signtx_group_bin_0078 = frame (4k)
frame_signtx_group_bin_0080 = frame (4k)
frame_signtx_group_bin_0081 = frame (4k)
frame_signtx_group_bin_0083 = frame (4k)
frame_signtx_group_bin_0084 = frame (4k)
frame_signtx_group_bin_0085 = frame (4k)
frame_signtx_group_bin_0086 = frame (4k)
frame_signtx_group_bin_0087 = frame (4k)
frame_signtx_group_bin_0088 = frame (4k)
frame_signtx_group_bin_0089 = frame (4k)
frame_signtx_group_bin_0090 = frame (4k)
frame_signtx_group_bin_0091 = frame (4k)
frame_signtx_group_bin_0092 = frame (4k)
frame_signtx_group_bin_0093 = frame (4k)
frame_signtx_group_bin_0094 = frame (4k)
frame_signtx_group_bin_0095 = frame (4k)
frame_signtx_group_bin_0096 = frame (4k)
frame_signtx_group_bin_0097 = frame (4k)
frame_signtx_group_bin_0098 = frame (4k)
frame_signtx_group_bin_0099 = frame (4k)
frame_signtx_group_bin_0100 = frame (4k)
frame_signtx_group_bin_0101 = frame (4k)
frame_signtx_group_bin_0102 = frame (4k)
frame_signtx_group_bin_0104 = frame (4k)
frame_signtx_group_bin_0105 = frame (4k)
frame_signtx_group_bin_0106 = frame (4k)
frame_signtx_group_bin_0107 = frame (4k)
frame_signtx_group_bin_0108 = frame (4k)
frame_signtx_group_bin_0109 = frame (4k)
frame_signtx_group_bin_0111 = frame (4k)
frame_signtx_group_bin_0112 = frame (4k)
frame_signtx_group_bin_0114 = frame (4k)
frame_signtx_group_bin_0115 = frame (4k)
frame_signtx_group_bin_0116 = frame (4k)
frame_signtx_group_bin_0117 = frame (4k)
frame_signtx_group_bin_0118 = frame (4k)
frame_signtx_group_bin_0119 = frame (4k)
frame_signtx_group_bin_0120 = frame (4k)
frame_signtx_group_bin_0121 = frame (4k)
frame_signtx_group_bin_0122 = frame (4k)
frame_signtx_group_bin_0123 = frame (4k)
frame_signtx_group_bin_0124 = frame (4k)
frame_signtx_group_bin_0125 = frame (4k)
frame_signtx_group_bin_0126 = frame (4k)
frame_signtx_group_bin_0127 = frame (4k)
frame_signtx_group_bin_0128 = frame (4k)
frame_signtx_group_bin_0129 = frame (4k)
frame_signtx_group_bin_0130 = frame (4k)
frame_signtx_group_bin_0131 = frame (4k)
frame_signtx_group_bin_0132 = frame (4k)
frame_signtx_group_bin_0133 = frame (4k)
frame_signtx_group_bin_0134 = frame (4k)
frame_signtx_group_bin_0136 = frame (4k)
frame_signtx_group_bin_0137 = frame (4k)
frame_signtx_group_bin_0138 = frame (4k)
frame_signtx_group_bin_0139 = frame (4k)
frame_signtx_group_bin_0140 = frame (4k)
frame_signtx_group_bin_0141 = frame (4k)
frame_signtx_group_bin_0142 = frame (4k)
frame_signtx_group_bin_0143 = frame (4k)
frame_signtx_group_bin_0144 = frame (4k)
frame_signtx_group_bin_0145 = frame (4k)
frame_signtx_group_bin_0146 = frame (4k)
frame_signtx_group_bin_0147 = frame (4k)
frame_signtx_group_bin_0148 = frame (4k)
frame_signtx_group_bin_0149 = frame (4k)
frame_signtx_group_bin_0151 = frame (4k)
frame_signtx_group_bin_0152 = frame (4k)
frame_signtx_group_bin_0153 = frame (4k)
frame_signtx_group_bin_0154 = frame (4k)
frame_signtx_group_bin_0155 = frame (4k)
frame_signtx_group_bin_0156 = frame (4k)
frame_signtx_group_bin_0158 = frame (4k)
frame_signtx_group_bin_0159 = frame (4k)
frame_signtx_group_bin_0160 = frame (4k)
frame_signtx_group_bin_0161 = frame (4k)
frame_signtx_group_bin_0162 = frame (4k)
frame_signtx_group_bin_0163 = frame (4k)
frame_signtx_group_bin_0164 = frame (4k)
frame_signtx_group_bin_0165 = frame (4k)
frame_signtx_group_bin_0166 = frame (4k)
frame_signtx_group_bin_0167 = frame (4k)
frame_signtx_group_bin_0168 = frame (4k)
frame_signtx_group_bin_0169 = frame (4k)
frame_signtx_group_bin_0170 = frame (4k)
frame_signtx_group_bin_0171 = frame (4k)
frame_signtx_group_bin_0172 = frame (4k)
frame_signtx_group_bin_0174 = frame (4k)
frame_signtx_group_bin_0175 = frame (4k)
frame_signtx_group_bin_0177 = frame (4k)
frame_signtx_group_bin_0178 = frame (4k)
frame_signtx_group_bin_0179 = frame (4k)
frame_signtx_group_bin_0180 = frame (4k)
frame_signtx_group_bin_0181 = frame (4k)
frame_signtx_group_bin_0182 = frame (4k)
frame_signtx_group_bin_0184 = frame (4k)
frame_signtx_group_bin_0185 = frame (4k)
frame_signtx_group_bin_0186 = frame (4k)
frame_signtx_group_bin_0187 = frame (4k)
frame_signtx_group_bin_0188 = frame (4k)
frame_signtx_group_bin_0189 = frame (4k)
frame_signtx_group_bin_0190 = frame (4k)
frame_signtx_group_bin_0191 = frame (4k)
frame_signtx_group_bin_0192 = frame (4k)
frame_signtx_group_bin_0193 = frame (4k)
frame_signtx_group_bin_0194 = frame (4k)
frame_signtx_group_bin_0195 = frame (4k)
frame_signtx_group_bin_0196 = frame (4k)
frame_signtx_group_bin_0197 = frame (4k)
frame_signtx_group_bin_0198 = frame (4k)
frame_signtx_group_bin_0199 = frame (4k)
frame_signtx_group_bin_0200 = frame (4k)
frame_signtx_group_bin_0201 = frame (4k)
frame_signtx_group_bin_0202 = frame (4k)
frame_signtx_group_bin_0203 = frame (4k)
frame_signtx_group_bin_0204 = frame (4k)
frame_signtx_group_bin_0205 = frame (4k)
frame_signtx_group_bin_0206 = frame (4k)
frame_signtx_group_bin_0207 = frame (4k)
frame_signtx_group_bin_0208 = frame (4k)
frame_signtx_group_bin_0209 = frame (4k)
frame_signtx_group_bin_0210 = frame (4k)
frame_signtx_group_bin_0211 = frame (4k)
frame_signtx_group_bin_0212 = frame (4k)
frame_signtx_group_bin_0213 = frame (4k)
frame_signtx_group_bin_0214 = frame (4k)
frame_signtx_group_bin_0215 = frame (4k)
frame_signtx_group_bin_0216 = frame (4k)
frame_signtx_group_bin_0217 = frame (4k)
frame_signtx_group_bin_0218 = frame (4k)
frame_signtx_group_bin_0219 = frame (4k)
frame_signtx_group_bin_0221 = frame (4k)
frame_signtx_group_bin_0222 = frame (4k)
frame_signtx_group_bin_0223 = frame (4k)
frame_signtx_group_bin_0224 = frame (4k)
frame_signtx_group_bin_0225 = frame (4k)
frame_signtx_group_bin_0226 = frame (4k)
frame_signtx_group_bin_0227 = frame (4k)
frame_signtx_group_bin_0229 = frame (4k)
frame_signtx_group_bin_0230 = frame (4k)
frame_signtx_group_bin_0231 = frame (4k)
frame_signtx_group_bin_0232 = frame (4k)
frame_signtx_group_bin_0233 = frame (4k)
frame_signtx_group_bin_0234 = frame (4k)
frame_signtx_group_bin_0235 = frame (4k)
frame_signtx_group_bin_0236 = frame (4k)
frame_signtx_group_bin_0237 = frame (4k)
frame_signtx_group_bin_0238 = frame (4k)
frame_signtx_group_bin_0239 = frame (4k)
frame_signtx_group_bin_0240 = frame (4k)
frame_signtx_group_bin_0241 = frame (4k)
frame_signtx_group_bin_0242 = frame (4k)
frame_signtx_group_bin_0243 = frame (4k)
frame_signtx_group_bin_0244 = frame (4k)
frame_signtx_group_bin_0245 = frame (4k)
frame_signtx_group_bin_0246 = frame (4k)
frame_signtx_group_bin_0247 = frame (4k)
frame_signtx_group_bin_0249 = frame (4k)
frame_signtx_group_bin_0250 = frame (4k)
frame_signtx_group_bin_0251 = frame (4k)
frame_signtx_group_bin_0252 = frame (4k)
frame_signtx_group_bin_0253 = frame (4k)
frame_signtx_group_bin_0254 = frame (4k)
frame_signtx_group_bin_0256 = frame (4k)
frame_signtx_group_bin_0257 = frame (4k)
frame_signtx_group_bin_0258 = frame (4k)
frame_signtx_group_bin_0259 = frame (4k)
frame_signtx_group_bin_0260 = frame (4k)
frame_signtx_group_bin_0261 = frame (4k)
frame_signtx_group_bin_0262 = frame (4k)
frame_signtx_group_bin_0263 = frame (4k)
frame_signtx_group_bin_0264 = frame (4k)
frame_signtx_group_bin_0265 = frame (4k)
frame_signtx_group_bin_0266 = frame (4k)
frame_signtx_group_bin_0267 = frame (4k)
frame_signtx_group_bin_0268 = frame (4k)
frame_signtx_group_bin_0269 = frame (4k)
frame_signtx_group_bin_0270 = frame (4k)
frame_signtx_group_bin_0271 = frame (4k)
frame_signtx_group_bin_0272 = frame (4k)
frame_signtx_group_bin_0273 = frame (4k)
frame_signtx_group_bin_0274 = frame (4k)
frame_signtx_group_bin_0275 = frame (4k)
frame_signtx_group_bin_0276 = frame (4k)
frame_signtx_group_bin_0277 = frame (4k)
frame_signtx_group_bin_0278 = frame (4k)
frame_signtx_group_bin_0279 = frame (4k)
frame_signtx_group_bin_0280 = frame (4k)
frame_signtx_group_bin_0281 = frame (4k)
frame_signtx_group_bin_0282 = frame (4k)
frame_signtx_group_bin_0283 = frame (4k)
frame_signtx_group_bin_0284 = frame (4k)
frame_signtx_group_bin_0285 = frame (4k)
frame_signtx_group_bin_0286 = frame (4k)
frame_signtx_group_bin_0287 = frame (4k)
frame_signtx_group_bin_0289 = frame (4k)
frame_signtx_group_bin_0290 = frame (4k)
frame_signtx_group_bin_0291 = frame (4k)
frame_signtx_group_bin_0292 = frame (4k)
frame_signtx_group_bin_0293 = frame (4k)
frame_signtx_group_bin_0294 = frame (4k)
frame_signtx_group_bin_0295 = frame (4k)
frame_signtx_group_bin_0296 = frame (4k)
frame_signtx_group_bin_0297 = frame (4k)
frame_signtx_group_bin_0298 = frame (4k)
frame_signtx_group_bin_0299 = frame (4k)
frame_signtx_group_bin_0300 = frame (4k)
frame_signtx_group_bin_0301 = frame (4k)
frame_signtx_group_bin_0302 = frame (4k)
frame_signtx_group_bin_0304 = frame (4k)
frame_signtx_group_bin_0305 = frame (4k)
frame_signtx_group_bin_0306 = frame (4k)
frame_signtx_group_bin_0307 = frame (4k)
frame_signtx_group_bin_0308 = frame (4k)
frame_signtx_group_bin_0309 = frame (4k)
frame_signtx_group_bin_0310 = frame (4k)
frame_signtx_group_bin_0311 = frame (4k)
frame_signtx_group_bin_0312 = frame (4k)
frame_signtx_group_bin_0313 = frame (4k)
frame_signtx_group_bin_0314 = frame (4k)
frame_signtx_group_bin_0315 = frame (4k)
frame_signtx_group_bin_0317 = frame (4k)
frame_signtx_group_bin_0319 = frame (4k)
frame_signtx_group_bin_0320 = frame (4k)
frame_signtx_group_bin_0321 = frame (4k)
frame_signtx_group_bin_0322 = frame (4k)
frame_signtx_group_bin_0323 = frame (4k)
frame_signtx_group_bin_0324 = frame (4k)
modchk_6_0_control_9_tcb = tcb (addr: 0x53cc00,ip: 0x406edd,sp: 0x52e000,elf: modchk_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [1],fault_ep: 0x00000002)
modchk_6_0_fault_handler_15_0000_tcb = tcb (addr: 0x542c00,ip: 0x406edd,sp: 0x53a000,elf: modchk_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [5])
modchk_6_modchk_iface_12_0000_tcb = tcb (addr: 0x53fc00,ip: 0x406edd,sp: 0x534000,elf: modchk_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [3],fault_ep: 0x00000004)
modchk_cnode = cnode (4 bits)
modchk_fault_ep = ep
modchk_frame__camkes_ipc_buffer_modchk_0_control = frame (4k)
modchk_frame__camkes_ipc_buffer_modchk_0_fault_handler_0000 = frame (4k)
modchk_frame__camkes_ipc_buffer_modchk_modchk_iface_0000 = frame (4k)
modchk_group_bin_pd = pml4
modchk_interface_init_ep = ep
modchk_post_init_ep = ep
modchk_pre_init_ep = ep
modtx_5_0_control_9_tcb = tcb (addr: 0x53bc00,ip: 0x40680e,sp: 0x52d000,elf: modtx_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [1],fault_ep: 0x00000002)
modtx_5_0_fault_handler_15_0000_tcb = tcb (addr: 0x541c00,ip: 0x40680e,sp: 0x539000,elf: modtx_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [5])
modtx_5_modtx_iface_11_0000_tcb = tcb (addr: 0x53ec00,ip: 0x40680e,sp: 0x533000,elf: modtx_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [3],fault_ep: 0x00000004)
modtx_cnode = cnode (4 bits)
modtx_fault_ep = ep
modtx_frame__camkes_ipc_buffer_modtx_0_control = frame (4k)
modtx_frame__camkes_ipc_buffer_modtx_0_fault_handler_0000 = frame (4k)
modtx_frame__camkes_ipc_buffer_modtx_modtx_iface_0000 = frame (4k)
modtx_group_bin_pd = pml4
modtx_interface_init_ep = ep
modtx_post_init_ep = ep
modtx_pre_init_ep = ep
pd_crypto_group_bin_0001 = pd
pd_modchk_group_bin_0001 = pd
pd_modtx_group_bin_0001 = pd
pd_signtx_group_bin_0001 = pd
pdpt_crypto_group_bin_0000 = pdpt
pdpt_modchk_group_bin_0000 = pdpt
pdpt_modtx_group_bin_0000 = pdpt
pdpt_signtx_group_bin_0000 = pdpt
pt_crypto_group_bin_0002 = pt
pt_modchk_group_bin_0002 = pt
pt_modtx_group_bin_0002 = pt
pt_signtx_group_bin_0002 = pt
signtx_6_0_control_9_tcb = tcb (addr: 0x53dc00,ip: 0x407bb4,sp: 0x52f000,elf: signtx_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [1],fault_ep: 0x00000002)
signtx_6_0_fault_handler_15_0000_tcb = tcb (addr: 0x543c00,ip: 0x407bb4,sp: 0x53b000,elf: signtx_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [5])
signtx_6_signtx_iface_12_0000_tcb = tcb (addr: 0x540c00,ip: 0x407bb4,sp: 0x535000,elf: signtx_group_bin,prio: 254,max_prio: 254,affinity: 0,init: [3],fault_ep: 0x00000004)
signtx_cnode = cnode (4 bits)
signtx_fault_ep = ep
signtx_frame__camkes_ipc_buffer_signtx_0_control = frame (4k)
signtx_frame__camkes_ipc_buffer_signtx_0_fault_handler_0000 = frame (4k)
signtx_frame__camkes_ipc_buffer_signtx_signtx_iface_0000 = frame (4k)
signtx_group_bin_pd = pml4
signtx_interface_init_ep = ep
signtx_post_init_ep = ep
signtx_pre_init_ep = ep
stack__camkes_stack_crypto_0_control_0_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_control_1_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_control_2_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_control_3_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_fault_handler_0000_0_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_fault_handler_0000_1_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_fault_handler_0000_2_crypto_obj = frame (4k)
stack__camkes_stack_crypto_0_fault_handler_0000_3_crypto_obj = frame (4k)
stack__camkes_stack_crypto_crypto_iface_0000_0_crypto_obj = frame (4k)
stack__camkes_stack_crypto_crypto_iface_0000_1_crypto_obj = frame (4k)
stack__camkes_stack_crypto_crypto_iface_0000_2_crypto_obj = frame (4k)
stack__camkes_stack_crypto_crypto_iface_0000_3_crypto_obj = frame (4k)
stack__camkes_stack_modchk_0_control_0_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_control_1_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_control_2_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_control_3_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_fault_handler_0000_0_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_fault_handler_0000_1_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_fault_handler_0000_2_modchk_obj = frame (4k)
stack__camkes_stack_modchk_0_fault_handler_0000_3_modchk_obj = frame (4k)
stack__camkes_stack_modchk_modchk_iface_0000_0_modchk_obj = frame (4k)
stack__camkes_stack_modchk_modchk_iface_0000_1_modchk_obj = frame (4k)
stack__camkes_stack_modchk_modchk_iface_0000_2_modchk_obj = frame (4k)
stack__camkes_stack_modchk_modchk_iface_0000_3_modchk_obj = frame (4k)
stack__camkes_stack_modtx_0_control_0_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_control_1_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_control_2_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_control_3_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_fault_handler_0000_0_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_fault_handler_0000_1_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_fault_handler_0000_2_modtx_obj = frame (4k)
stack__camkes_stack_modtx_0_fault_handler_0000_3_modtx_obj = frame (4k)
stack__camkes_stack_modtx_modtx_iface_0000_0_modtx_obj = frame (4k)
stack__camkes_stack_modtx_modtx_iface_0000_1_modtx_obj = frame (4k)
stack__camkes_stack_modtx_modtx_iface_0000_2_modtx_obj = frame (4k)
stack__camkes_stack_modtx_modtx_iface_0000_3_modtx_obj = frame (4k)
stack__camkes_stack_signtx_0_control_0_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_control_1_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_control_2_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_control_3_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_fault_handler_0000_0_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_fault_handler_0000_1_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_fault_handler_0000_2_signtx_obj = frame (4k)
stack__camkes_stack_signtx_0_fault_handler_0000_3_signtx_obj = frame (4k)
stack__camkes_stack_signtx_signtx_iface_0000_0_signtx_obj = frame (4k)
stack__camkes_stack_signtx_signtx_iface_0000_1_signtx_obj = frame (4k)
stack__camkes_stack_signtx_signtx_iface_0000_2_signtx_obj = frame (4k)
stack__camkes_stack_signtx_signtx_iface_0000_3_signtx_obj = frame (4k)
}

caps {
crypto_6_0_control_9_tcb {
cspace: crypto_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: crypto_frame__camkes_ipc_buffer_crypto_0_control (RW)
vspace: crypto_group_bin_pd
}
crypto_6_0_fault_handler_15_0000_tcb {
cspace: crypto_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: crypto_frame__camkes_ipc_buffer_crypto_0_fault_handler_0000 (RW)
vspace: crypto_group_bin_pd
}
crypto_6_crypto_iface_12_0000_tcb {
cspace: crypto_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: crypto_frame__camkes_ipc_buffer_crypto_crypto_iface_0000 (RW)
vspace: crypto_group_bin_pd
}
crypto_cnode {
0x1: crypto_6_0_control_9_tcb
0x2: crypto_fault_ep (RWX, badge: 1)
0x3: crypto_6_crypto_iface_12_0000_tcb
0x4: crypto_fault_ep (RWX, badge: 3)
0x5: crypto_6_0_fault_handler_15_0000_tcb
0x6: crypto_fault_ep (RWX)
0x7: crypto_pre_init_ep (RW)
0x8: crypto_interface_init_ep (RW)
0x9: crypto_post_init_ep (RW)
0xa: conn2.conn5_ep (RW)
0xb: crypto_cnode (guard: 0, guard_size: 60)
0xd: conn3.conn7_ep (WX, badge: 1)
0xe: conn4.conn8_ep (WX, badge: 1)
}
crypto_group_bin_pd {
0x0: pdpt_crypto_group_bin_0000
}
modchk_6_0_control_9_tcb {
cspace: modchk_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: modchk_frame__camkes_ipc_buffer_modchk_0_control (RW)
vspace: modchk_group_bin_pd
}
modchk_6_0_fault_handler_15_0000_tcb {
cspace: modchk_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: modchk_frame__camkes_ipc_buffer_modchk_0_fault_handler_0000 (RW)
vspace: modchk_group_bin_pd
}
modchk_6_modchk_iface_12_0000_tcb {
cspace: modchk_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: modchk_frame__camkes_ipc_buffer_modchk_modchk_iface_0000 (RW)
vspace: modchk_group_bin_pd
}
modchk_cnode {
0x1: modchk_6_0_control_9_tcb
0x2: modchk_fault_ep (RWX, badge: 1)
0x3: modchk_6_modchk_iface_12_0000_tcb
0x4: modchk_fault_ep (RWX, badge: 3)
0x5: modchk_6_0_fault_handler_15_0000_tcb
0x6: modchk_fault_ep (RWX)
0x7: modchk_pre_init_ep (RW)
0x8: modchk_interface_init_ep (RW)
0x9: modchk_post_init_ep (RW)
0xa: conn1.conn6_ep (RW)
0xb: modchk_cnode (guard: 0, guard_size: 60)
0xd: conn3.conn7_ep (WX, badge: 2)
0xe: conn4.conn8_ep (WX, badge: 2)
}
modchk_group_bin_pd {
0x0: pdpt_modchk_group_bin_0000
}
modtx_5_0_control_9_tcb {
cspace: modtx_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: modtx_frame__camkes_ipc_buffer_modtx_0_control (RW)
vspace: modtx_group_bin_pd
}
modtx_5_0_fault_handler_15_0000_tcb {
cspace: modtx_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: modtx_frame__camkes_ipc_buffer_modtx_0_fault_handler_0000 (RW)
vspace: modtx_group_bin_pd
}
modtx_5_modtx_iface_11_0000_tcb {
cspace: modtx_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: modtx_frame__camkes_ipc_buffer_modtx_modtx_iface_0000 (RW)
vspace: modtx_group_bin_pd
}
modtx_cnode {
0x1: modtx_5_0_control_9_tcb
0x2: modtx_fault_ep (RWX, badge: 1)
0x3: modtx_5_modtx_iface_11_0000_tcb
0x4: modtx_fault_ep (RWX, badge: 3)
0x5: modtx_5_0_fault_handler_15_0000_tcb
0x6: modtx_fault_ep (RWX)
0x7: modtx_pre_init_ep (RW)
0x8: modtx_interface_init_ep (RW)
0x9: modtx_post_init_ep (RW)
0xa: conn2.conn5_ep (WX, badge: 1)
0xb: conn1.conn6_ep (WX, badge: 1)
0xc: conn3.conn7_ep (RW)
0xd: modtx_cnode (guard: 0, guard_size: 60)
}
modtx_group_bin_pd {
0x0: pdpt_modtx_group_bin_0000
}
pd_crypto_group_bin_0001 {
0x2: pt_crypto_group_bin_0002
}
pd_modchk_group_bin_0001 {
0x2: pt_modchk_group_bin_0002
}
pd_modtx_group_bin_0001 {
0x2: pt_modtx_group_bin_0002
}
pd_signtx_group_bin_0001 {
0x2: pt_signtx_group_bin_0002
}
pdpt_crypto_group_bin_0000 {
0x0: pd_crypto_group_bin_0001
}
pdpt_modchk_group_bin_0000 {
0x0: pd_modchk_group_bin_0001
}
pdpt_modtx_group_bin_0000 {
0x0: pd_modtx_group_bin_0001
}
pdpt_signtx_group_bin_0000 {
0x0: pd_signtx_group_bin_0001
}
pt_crypto_group_bin_0002 {
0x0: frame_crypto_group_bin_0000 (RX)
0x100: frame_crypto_group_bin_0030 (RW)
0x101: frame_crypto_group_bin_0180 (RW)
0x102: frame_crypto_group_bin_0233 (RW)
0x103: frame_crypto_group_bin_0160 (RW)
0x104: frame_crypto_group_bin_0285 (RW)
0x105: frame_crypto_group_bin_0107 (RW)
0x106: frame_crypto_group_bin_0252 (RW)
0x107: frame_crypto_group_bin_0298 (RW)
0x108: frame_crypto_group_bin_0304 (RW)
0x109: frame_crypto_group_bin_0072 (RW)
0x10: frame_crypto_group_bin_0060 (RX)
0x10a: frame_crypto_group_bin_0167 (RW)
0x10b: frame_crypto_group_bin_0261 (RW)
0x10c: frame_crypto_group_bin_0027 (RW)
0x10d: frame_crypto_group_bin_0125 (RW)
0x10e: frame_crypto_group_bin_0217 (RW)
0x10f: frame_crypto_group_bin_0311 (RW)
0x110: frame_crypto_group_bin_0080 (RW)
0x111: frame_crypto_group_bin_0177 (RW)
0x112: frame_crypto_group_bin_0111 (RW)
0x113: frame_crypto_group_bin_0037 (RW)
0x114: frame_crypto_group_bin_0133 (RW)
0x115: frame_crypto_group_bin_0224 (RW)
0x116: frame_crypto_group_bin_0319 (RW)
0x117: frame_crypto_group_bin_0089 (RW)
0x118: frame_crypto_group_bin_0265 (RW)
0x119: frame_crypto_group_bin_0086 (RW)
0x11: frame_crypto_group_bin_0146 (RX)
0x11a: frame_crypto_group_bin_0174 (RW)
0x11b: frame_crypto_group_bin_0098 (RW)
0x11c: frame_crypto_group_bin_0195 (RW)
0x11d: frame_crypto_group_bin_0014 (RW)
0x11e: frame_crypto_group_bin_0161 (RW)
0x11f: frame_crypto_group_bin_0192 (RW)
0x120: frame_crypto_group_bin_0284 (RW)
0x121: frame_crypto_group_bin_0270 (RW)
0x122: frame_crypto_group_bin_0237 (RW)
0x123: frame_crypto_group_bin_0024 (RW)
0x124: frame_crypto_group_bin_0054 (RW)
0x125: frame_crypto_group_bin_0201 (RW)
0x126: frame_crypto_group_bin_0019 (RW)
0x127: frame_crypto_group_bin_0293 (RW)
0x128: frame_crypto_group_bin_0260 (RW)
0x129: frame_crypto_group_bin_0009 (RW)
0x12: frame_crypto_group_bin_0227 (RX)
0x12b: stack__camkes_stack_crypto_0_control_0_crypto_obj (RW)
0x12c: stack__camkes_stack_crypto_0_control_1_crypto_obj (RW)
0x12d: stack__camkes_stack_crypto_0_control_2_crypto_obj (RW)
0x12e: stack__camkes_stack_crypto_0_control_3_crypto_obj (RW)
0x131: stack__camkes_stack_crypto_crypto_iface_0000_0_crypto_obj (RW)
0x132: stack__camkes_stack_crypto_crypto_iface_0000_1_crypto_obj (RW)
0x133: stack__camkes_stack_crypto_crypto_iface_0000_2_crypto_obj (RW)
0x134: stack__camkes_stack_crypto_crypto_iface_0000_3_crypto_obj (RW)
0x137: stack__camkes_stack_crypto_0_fault_handler_0000_0_crypto_obj (RW)
0x138: stack__camkes_stack_crypto_0_fault_handler_0000_1_crypto_obj (RW)
0x139: stack__camkes_stack_crypto_0_fault_handler_0000_2_crypto_obj (RW)
0x13: frame_crypto_group_bin_0312 (RX)
0x13a: stack__camkes_stack_crypto_0_fault_handler_0000_3_crypto_obj (RW)
0x13d: crypto_frame__camkes_ipc_buffer_crypto_0_control (RW)
0x140: crypto_frame__camkes_ipc_buffer_crypto_crypto_iface_0000 (RW)
0x143: crypto_frame__camkes_ipc_buffer_crypto_0_fault_handler_0000 (RW)
0x14: frame_crypto_group_bin_0071 (RX)
0x15: frame_crypto_group_bin_0156 (RX)
0x16: frame_crypto_group_bin_0239 (RX)
0x17: frame_crypto_group_bin_0322 (RX)
0x18: frame_crypto_group_bin_0081 (RX)
0x19: frame_crypto_group_bin_0087 (RX)
0x1: frame_crypto_group_bin_0001 (RX)
0x1a: frame_crypto_group_bin_0250 (RX)
0x1b: frame_crypto_group_bin_0249 (RX)
0x1c: frame_crypto_group_bin_0004 (RX)
0x1d: frame_crypto_group_bin_0178 (RX)
0x1e: frame_crypto_group_bin_0259 (RX)
0x1f: frame_crypto_group_bin_0017 (RX)
0x20: frame_crypto_group_bin_0102 (RX)
0x21: frame_crypto_group_bin_0187 (RX)
0x22: frame_crypto_group_bin_0268 (RX)
0x23: frame_crypto_group_bin_0026 (RX)
0x24: frame_crypto_group_bin_0115 (RX)
0x25: frame_crypto_group_bin_0197 (RX)
0x26: frame_crypto_group_bin_0278 (RW)
0x27: frame_crypto_group_bin_0038 (RW)
0x28: frame_crypto_group_bin_0124 (RW)
0x29: frame_crypto_group_bin_0207 (RW)
0x2: frame_crypto_group_bin_0190 (RX)
0x2a: frame_crypto_group_bin_0290 (RW)
0x2b: frame_crypto_group_bin_0047 (RW)
0x2c: frame_crypto_group_bin_0134 (RW)
0x2d: frame_crypto_group_bin_0216 (RW)
0x2e: frame_crypto_group_bin_0300 (RW)
0x2f: frame_crypto_group_bin_0058 (RW)
0x30: frame_crypto_group_bin_0144 (RW)
0x31: frame_crypto_group_bin_0225 (RW)
0x32: frame_crypto_group_bin_0310 (RW)
0x33: frame_crypto_group_bin_0068 (RW)
0x34: frame_crypto_group_bin_0154 (RW)
0x35: frame_crypto_group_bin_0235 (RW)
0x36: frame_crypto_group_bin_0320 (RW)
0x37: frame_crypto_group_bin_0078 (RW)
0x38: frame_crypto_group_bin_0164 (RW)
0x39: frame_crypto_group_bin_0247 (RW)
0x3: frame_crypto_group_bin_0271 (RX)
0x3a: frame_crypto_group_bin_0168 (RW)
0x3b: frame_crypto_group_bin_0090 (RW)
0x3c: frame_crypto_group_bin_0175 (RW)
0x3d: frame_crypto_group_bin_0257 (RW)
0x3e: frame_crypto_group_bin_0015 (RW)
0x3f: frame_crypto_group_bin_0099 (RW)
0x40: frame_crypto_group_bin_0185 (RW)
0x41: frame_crypto_group_bin_0266 (RW)
0x42: frame_crypto_group_bin_0023 (RW)
0x43: frame_crypto_group_bin_0112 (RW)
0x44: frame_crypto_group_bin_0194 (RW)
0x45: frame_crypto_group_bin_0276 (RW)
0x46: frame_crypto_group_bin_0035 (RW)
0x47: frame_crypto_group_bin_0122 (RW)
0x48: frame_crypto_group_bin_0204 (RW)
0x49: frame_crypto_group_bin_0286 (RW)
0x4: frame_crypto_group_bin_0028 (RX)
0x4a: frame_crypto_group_bin_0045 (RW)
0x4b: frame_crypto_group_bin_0131 (RW)
0x4c: frame_crypto_group_bin_0213 (RW)
0x4d: frame_crypto_group_bin_0297 (RW)
0x4e: frame_crypto_group_bin_0055 (RW)
0x4f: frame_crypto_group_bin_0142 (RW)
0x50: frame_crypto_group_bin_0223 (RW)
0x51: frame_crypto_group_bin_0307 (RW)
0x52: frame_crypto_group_bin_0065 (RW)
0x53: frame_crypto_group_bin_0151 (RW)
0x54: frame_crypto_group_bin_0232 (RW)
0x55: frame_crypto_group_bin_0317 (RW)
0x56: frame_crypto_group_bin_0075 (RW)
0x57: frame_crypto_group_bin_0162 (RW)
0x58: frame_crypto_group_bin_0244 (RW)
0x59: frame_crypto_group_bin_0002 (RW)
0x5: frame_crypto_group_bin_0118 (RX)
0x5a: frame_crypto_group_bin_0088 (RW)
0x5b: frame_crypto_group_bin_0171 (RW)
0x5c: frame_crypto_group_bin_0256 (RW)
0x5d: frame_crypto_group_bin_0013 (RW)
0x5e: frame_crypto_group_bin_0097 (RW)
0x5f: frame_crypto_group_bin_0184 (RW)
0x60: frame_crypto_group_bin_0264 (RW)
0x61: frame_crypto_group_bin_0022 (RW)
0x62: frame_crypto_group_bin_0108 (RW)
0x63: frame_crypto_group_bin_0193 (RW)
0x64: frame_crypto_group_bin_0273 (RW)
0x65: frame_crypto_group_bin_0031 (RW)
0x66: frame_crypto_group_bin_0120 (RW)
0x67: frame_crypto_group_bin_0202 (RW)
0x68: frame_crypto_group_bin_0283 (RW)
0x69: frame_crypto_group_bin_0043 (RW)
0x6: frame_crypto_group_bin_0199 (RX)
0x6a: frame_crypto_group_bin_0128 (RW)
0x6b: frame_crypto_group_bin_0211 (RW)
0x6c: frame_crypto_group_bin_0295 (RW)
0x6d: frame_crypto_group_bin_0052 (RW)
0x6e: frame_crypto_group_bin_0140 (RW)
0x6f: frame_crypto_group_bin_0221 (RW)
0x70: frame_crypto_group_bin_0305 (RW)
0x71: frame_crypto_group_bin_0062 (RW)
0x72: frame_crypto_group_bin_0148 (RW)
0x73: frame_crypto_group_bin_0230 (RW)
0x74: frame_crypto_group_bin_0314 (RW)
0x75: frame_crypto_group_bin_0073 (RW)
0x76: frame_crypto_group_bin_0159 (RW)
0x77: frame_crypto_group_bin_0241 (RW)
0x78: frame_crypto_group_bin_0324 (RW)
0x79: frame_crypto_group_bin_0084 (RW)
0x7: frame_crypto_group_bin_0281 (RX)
0x7a: frame_crypto_group_bin_0169 (RW)
0x7b: frame_crypto_group_bin_0253 (RW)
0x7c: frame_crypto_group_bin_0011 (RW)
0x7d: frame_crypto_group_bin_0095 (RW)
0x7e: frame_crypto_group_bin_0181 (RW)
0x7f: frame_crypto_group_bin_0262 (RW)
0x80: frame_crypto_group_bin_0020 (RW)
0x81: frame_crypto_group_bin_0105 (RW)
0x82: frame_crypto_group_bin_0053 (RW)
0x83: frame_crypto_group_bin_0149 (RW)
0x84: frame_crypto_group_bin_0242 (RW)
0x85: frame_crypto_group_bin_0012 (RW)
0x86: frame_crypto_group_bin_0106 (RW)
0x87: frame_crypto_group_bin_0200 (RW)
0x88: frame_crypto_group_bin_0294 (RW)
0x89: frame_crypto_group_bin_0061 (RW)
0x8: frame_crypto_group_bin_0041 (RX)
0x8a: frame_crypto_group_bin_0158 (RW)
0x8b: frame_crypto_group_bin_0251 (RW)
0x8c: frame_crypto_group_bin_0018 (RW)
0x8d: frame_crypto_group_bin_0117 (RW)
0x8e: frame_crypto_group_bin_0208 (RW)
0x8f: frame_crypto_group_bin_0301 (RW)
0x90: frame_crypto_group_bin_0070 (RW)
0x91: frame_crypto_group_bin_0165 (RW)
0x92: frame_crypto_group_bin_0258 (RW)
0x93: frame_crypto_group_bin_0025 (RW)
0x94: frame_crypto_group_bin_0123 (RW)
0x95: frame_crypto_group_bin_0215 (RW)
0x96: frame_crypto_group_bin_0309 (RW)
0x97: frame_crypto_group_bin_0077 (RW)
0x98: frame_crypto_group_bin_0214 (RW)
0x99: frame_crypto_group_bin_0166 (RW)
0x9: frame_crypto_group_bin_0126 (RX)
0x9a: frame_crypto_group_bin_0182 (RW)
0x9b: frame_crypto_group_bin_0008 (RW)
0x9c: frame_crypto_group_bin_0092 (RW)
0x9d: frame_crypto_group_bin_0287 (RW)
0x9e: frame_crypto_group_bin_0109 (RW)
0x9f: frame_crypto_group_bin_0254 (RW)
0xa0: frame_crypto_group_bin_0274 (RW)
0xa1: frame_crypto_group_bin_0044 (RW)
0xa2: frame_crypto_group_bin_0141 (RW)
0xa3: frame_crypto_group_bin_0231 (RW)
0xa4: frame_crypto_group_bin_0003 (RW)
0xa5: frame_crypto_group_bin_0096 (RW)
0xa6: frame_crypto_group_bin_0191 (RW)
0xa7: frame_crypto_group_bin_0282 (RW)
0xa8: frame_crypto_group_bin_0051 (RW)
0xa9: frame_crypto_group_bin_0147 (RW)
0xa: frame_crypto_group_bin_0209 (RX)
0xaa: frame_crypto_group_bin_0240 (RW)
0xab: frame_crypto_group_bin_0010 (RW)
0xac: frame_crypto_group_bin_0104 (RW)
0xad: frame_crypto_group_bin_0198 (RW)
0xae: frame_crypto_group_bin_0291 (RW)
0xaf: frame_crypto_group_bin_0059 (RW)
0xb0: frame_crypto_group_bin_0155 (RW)
0xb1: frame_crypto_group_bin_0029 (RW)
0xb2: frame_crypto_group_bin_0016 (RW)
0xb3: frame_crypto_group_bin_0114 (RW)
0xb4: frame_crypto_group_bin_0206 (RW)
0xb5: frame_crypto_group_bin_0299 (RW)
0xb6: frame_crypto_group_bin_0067 (RW)
0xb7: frame_crypto_group_bin_0163 (RW)
0xb8: frame_crypto_group_bin_0308 (RW)
0xb9: frame_crypto_group_bin_0129 (RW)
0xb: frame_crypto_group_bin_0292 (RX)
0xba: frame_crypto_group_bin_0005 (RW)
0xbb: frame_crypto_group_bin_0093 (RW)
0xbc: frame_crypto_group_bin_0236 (RW)
0xbd: frame_crypto_group_bin_0056 (RW)
0xbe: frame_crypto_group_bin_0203 (RW)
0xbf: frame_crypto_group_bin_0021 (RW)
0xc0: frame_crypto_group_bin_0032 (RW)
0xc1: frame_crypto_group_bin_0313 (RW)
0xc2: frame_crypto_group_bin_0222 (RW)
0xc3: frame_crypto_group_bin_0315 (RW)
0xc4: frame_crypto_group_bin_0085 (RW)
0xc5: frame_crypto_group_bin_0243 (RW)
0xc6: frame_crypto_group_bin_0272 (RW)
0xc7: frame_crypto_group_bin_0042 (RW)
0xc8: frame_crypto_group_bin_0139 (RW)
0xc9: frame_crypto_group_bin_0229 (RW)
0xc: frame_crypto_group_bin_0049 (RX)
0xca: frame_crypto_group_bin_0323 (RW)
0xcb: frame_crypto_group_bin_0094 (RW)
0xcc: frame_crypto_group_bin_0189 (RW)
0xcd: frame_crypto_group_bin_0280 (RW)
0xce: frame_crypto_group_bin_0048 (RW)
0xcf: frame_crypto_group_bin_0145 (RW)
0xd0: frame_crypto_group_bin_0238 (RW)
0xd1: frame_crypto_group_bin_0007 (RW)
0xd2: frame_crypto_group_bin_0101 (RW)
0xd3: frame_crypto_group_bin_0196 (RW)
0xd4: frame_crypto_group_bin_0289 (RW)
0xd5: frame_crypto_group_bin_0057 (RW)
0xd6: frame_crypto_group_bin_0153 (RW)
0xd7: frame_crypto_group_bin_0246 (RW)
0xd8: frame_crypto_group_bin_0076 (RW)
0xd9: frame_crypto_group_bin_0132 (RW)
0xd: frame_crypto_group_bin_0137 (RX)
0xda: frame_crypto_group_bin_0205 (RW)
0xdb: frame_crypto_group_bin_0188 (RW)
0xdc: frame_crypto_group_bin_0006 (RW)
0xdd: frame_crypto_group_bin_0152 (RW)
0xde: frame_crypto_group_bin_0296 (RW)
0xdf: frame_crypto_group_bin_0119 (RW)
0xe0: frame_crypto_group_bin_0121 (RW)
0xe1: frame_crypto_group_bin_0212 (RW)
0xe2: frame_crypto_group_bin_0306 (RW)
0xe3: frame_crypto_group_bin_0074 (RW)
0xe4: frame_crypto_group_bin_0170 (RW)
0xe5: frame_crypto_group_bin_0263 (RW)
0xe6: frame_crypto_group_bin_0130 (RW)
0xe7: frame_crypto_group_bin_0127 (RW)
0xe8: frame_crypto_group_bin_0219 (RW)
0xe9: frame_crypto_group_bin_0267 (RW)
0xe: frame_crypto_group_bin_0218 (RX)
0xea: frame_crypto_group_bin_0083 (RW)
0xeb: frame_crypto_group_bin_0179 (RW)
0xec: frame_crypto_group_bin_0269 (RW)
0xed: frame_crypto_group_bin_0039 (RW)
0xee: frame_crypto_group_bin_0136 (RW)
0xef: frame_crypto_group_bin_0226 (RW)
0xf0: frame_crypto_group_bin_0321 (RW)
0xf1: frame_crypto_group_bin_0091 (RW)
0xf2: frame_crypto_group_bin_0186 (RW)
0xf3: frame_crypto_group_bin_0277 (RW)
0xf4: frame_crypto_group_bin_0046 (RW)
0xf5: frame_crypto_group_bin_0143 (RW)
0xf6: frame_crypto_group_bin_0234 (RW)
0xf7: frame_crypto_group_bin_0116 (RW)
0xf8: frame_crypto_group_bin_0172 (RW)
0xf9: frame_crypto_group_bin_0275 (RW)
0xf: frame_crypto_group_bin_0302 (RX)
0xfa: frame_crypto_group_bin_0138 (RW)
0xfb: frame_crypto_group_bin_0279 (RW)
0xfc: frame_crypto_group_bin_0100 (RW)
0xfd: frame_crypto_group_bin_0245 (RW)
0xfe: frame_crypto_group_bin_0063 (RW)
0xff: frame_crypto_group_bin_0210 (RW)
}
pt_modchk_group_bin_0002 {
0x0: frame_modchk_group_bin_0000 (RX)
0x100: frame_modchk_group_bin_0030 (RW)
0x101: frame_modchk_group_bin_0179 (RW)
0x102: frame_modchk_group_bin_0232 (RW)
0x103: frame_modchk_group_bin_0159 (RW)
0x104: frame_modchk_group_bin_0284 (RW)
0x105: frame_modchk_group_bin_0107 (RW)
0x106: frame_modchk_group_bin_0251 (RW)
0x107: frame_modchk_group_bin_0297 (RW)
0x108: frame_modchk_group_bin_0303 (RW)
0x109: frame_modchk_group_bin_0072 (RW)
0x10: frame_modchk_group_bin_0060 (RX)
0x10a: frame_modchk_group_bin_0166 (RW)
0x10b: frame_modchk_group_bin_0260 (RW)
0x10c: frame_modchk_group_bin_0027 (RW)
0x10d: frame_modchk_group_bin_0125 (RW)
0x10e: frame_modchk_group_bin_0216 (RW)
0x10f: frame_modchk_group_bin_0310 (RW)
0x110: frame_modchk_group_bin_0080 (RW)
0x111: frame_modchk_group_bin_0176 (RW)
0x112: frame_modchk_group_bin_0111 (RW)
0x113: frame_modchk_group_bin_0037 (RW)
0x114: frame_modchk_group_bin_0133 (RW)
0x115: frame_modchk_group_bin_0223 (RW)
0x116: frame_modchk_group_bin_0318 (RW)
0x117: frame_modchk_group_bin_0089 (RW)
0x118: frame_modchk_group_bin_0264 (RW)
0x119: frame_modchk_group_bin_0086 (RW)
0x11: frame_modchk_group_bin_0146 (RX)
0x11a: frame_modchk_group_bin_0173 (RW)
0x11b: frame_modchk_group_bin_0098 (RW)
0x11c: frame_modchk_group_bin_0194 (RW)
0x11d: frame_modchk_group_bin_0014 (RW)
0x11e: frame_modchk_group_bin_0160 (RW)
0x11f: frame_modchk_group_bin_0191 (RW)
0x120: frame_modchk_group_bin_0283 (RW)
0x121: frame_modchk_group_bin_0269 (RW)
0x122: frame_modchk_group_bin_0236 (RW)
0x123: frame_modchk_group_bin_0024 (RW)
0x124: frame_modchk_group_bin_0054 (RW)
0x125: frame_modchk_group_bin_0200 (RW)
0x126: frame_modchk_group_bin_0019 (RW)
0x127: frame_modchk_group_bin_0292 (RW)
0x128: frame_modchk_group_bin_0259 (RW)
0x12: frame_modchk_group_bin_0226 (RX)
0x12a: stack__camkes_stack_modchk_0_control_0_modchk_obj (RW)
0x12b: stack__camkes_stack_modchk_0_control_1_modchk_obj (RW)
0x12c: stack__camkes_stack_modchk_0_control_2_modchk_obj (RW)
0x12d: stack__camkes_stack_modchk_0_control_3_modchk_obj (RW)
0x130: stack__camkes_stack_modchk_modchk_iface_0000_0_modchk_obj (RW)
0x131: stack__camkes_stack_modchk_modchk_iface_0000_1_modchk_obj (RW)
0x132: stack__camkes_stack_modchk_modchk_iface_0000_2_modchk_obj (RW)
0x133: stack__camkes_stack_modchk_modchk_iface_0000_3_modchk_obj (RW)
0x136: stack__camkes_stack_modchk_0_fault_handler_0000_0_modchk_obj (RW)
0x137: stack__camkes_stack_modchk_0_fault_handler_0000_1_modchk_obj (RW)
0x138: stack__camkes_stack_modchk_0_fault_handler_0000_2_modchk_obj (RW)
0x139: stack__camkes_stack_modchk_0_fault_handler_0000_3_modchk_obj (RW)
0x13: frame_modchk_group_bin_0311 (RX)
0x13c: modchk_frame__camkes_ipc_buffer_modchk_0_control (RW)
0x13f: modchk_frame__camkes_ipc_buffer_modchk_modchk_iface_0000 (RW)
0x142: modchk_frame__camkes_ipc_buffer_modchk_0_fault_handler_0000 (RW)
0x14: frame_modchk_group_bin_0071 (RX)
0x15: frame_modchk_group_bin_0155 (RX)
0x16: frame_modchk_group_bin_0238 (RX)
0x17: frame_modchk_group_bin_0321 (RX)
0x18: frame_modchk_group_bin_0081 (RX)
0x19: frame_modchk_group_bin_0087 (RX)
0x1: frame_modchk_group_bin_0001 (RX)
0x1a: frame_modchk_group_bin_0249 (RX)
0x1b: frame_modchk_group_bin_0248 (RX)
0x1c: frame_modchk_group_bin_0004 (RX)
0x1d: frame_modchk_group_bin_0177 (RX)
0x1e: frame_modchk_group_bin_0258 (RX)
0x1f: frame_modchk_group_bin_0017 (RX)
0x20: frame_modchk_group_bin_0102 (RX)
0x21: frame_modchk_group_bin_0186 (RX)
0x22: frame_modchk_group_bin_0267 (RX)
0x23: frame_modchk_group_bin_0026 (RX)
0x24: frame_modchk_group_bin_0115 (RX)
0x25: frame_modchk_group_bin_0196 (RW)
0x26: frame_modchk_group_bin_0277 (RW)
0x27: frame_modchk_group_bin_0038 (RW)
0x28: frame_modchk_group_bin_0124 (RW)
0x29: frame_modchk_group_bin_0206 (RW)
0x2: frame_modchk_group_bin_0189 (RX)
0x2a: frame_modchk_group_bin_0289 (RW)
0x2b: frame_modchk_group_bin_0047 (RW)
0x2c: frame_modchk_group_bin_0134 (RW)
0x2d: frame_modchk_group_bin_0215 (RW)
0x2e: frame_modchk_group_bin_0299 (RW)
0x2f: frame_modchk_group_bin_0058 (RW)
0x30: frame_modchk_group_bin_0144 (RW)
0x31: frame_modchk_group_bin_0224 (RW)
0x32: frame_modchk_group_bin_0309 (RW)
0x33: frame_modchk_group_bin_0068 (RW)
0x34: frame_modchk_group_bin_0153 (RW)
0x35: frame_modchk_group_bin_0234 (RW)
0x36: frame_modchk_group_bin_0319 (RW)
0x37: frame_modchk_group_bin_0078 (RW)
0x38: frame_modchk_group_bin_0163 (RW)
0x39: frame_modchk_group_bin_0246 (RW)
0x3: frame_modchk_group_bin_0270 (RX)
0x3a: frame_modchk_group_bin_0167 (RW)
0x3b: frame_modchk_group_bin_0090 (RW)
0x3c: frame_modchk_group_bin_0174 (RW)
0x3d: frame_modchk_group_bin_0256 (RW)
0x3e: frame_modchk_group_bin_0015 (RW)
0x3f: frame_modchk_group_bin_0099 (RW)
0x40: frame_modchk_group_bin_0184 (RW)
0x41: frame_modchk_group_bin_0265 (RW)
0x42: frame_modchk_group_bin_0023 (RW)
0x43: frame_modchk_group_bin_0112 (RW)
0x44: frame_modchk_group_bin_0193 (RW)
0x45: frame_modchk_group_bin_0275 (RW)
0x46: frame_modchk_group_bin_0035 (RW)
0x47: frame_modchk_group_bin_0122 (RW)
0x48: frame_modchk_group_bin_0203 (RW)
0x49: frame_modchk_group_bin_0285 (RW)
0x4: frame_modchk_group_bin_0028 (RX)
0x4a: frame_modchk_group_bin_0045 (RW)
0x4b: frame_modchk_group_bin_0131 (RW)
0x4c: frame_modchk_group_bin_0212 (RW)
0x4d: frame_modchk_group_bin_0296 (RW)
0x4e: frame_modchk_group_bin_0055 (RW)
0x4f: frame_modchk_group_bin_0142 (RW)
0x50: frame_modchk_group_bin_0222 (RW)
0x51: frame_modchk_group_bin_0306 (RW)
0x52: frame_modchk_group_bin_0065 (RW)
0x53: frame_modchk_group_bin_0150 (RW)
0x54: frame_modchk_group_bin_0231 (RW)
0x55: frame_modchk_group_bin_0316 (RW)
0x56: frame_modchk_group_bin_0075 (RW)
0x57: frame_modchk_group_bin_0161 (RW)
0x58: frame_modchk_group_bin_0243 (RW)
0x59: frame_modchk_group_bin_0002 (RW)
0x5: frame_modchk_group_bin_0118 (RX)
0x5a: frame_modchk_group_bin_0088 (RW)
0x5b: frame_modchk_group_bin_0170 (RW)
0x5c: frame_modchk_group_bin_0255 (RW)
0x5d: frame_modchk_group_bin_0013 (RW)
0x5e: frame_modchk_group_bin_0097 (RW)
0x5f: frame_modchk_group_bin_0183 (RW)
0x60: frame_modchk_group_bin_0263 (RW)
0x61: frame_modchk_group_bin_0022 (RW)
0x62: frame_modchk_group_bin_0108 (RW)
0x63: frame_modchk_group_bin_0192 (RW)
0x64: frame_modchk_group_bin_0272 (RW)
0x65: frame_modchk_group_bin_0031 (RW)
0x66: frame_modchk_group_bin_0120 (RW)
0x67: frame_modchk_group_bin_0201 (RW)
0x68: frame_modchk_group_bin_0282 (RW)
0x69: frame_modchk_group_bin_0043 (RW)
0x6: frame_modchk_group_bin_0198 (RX)
0x6a: frame_modchk_group_bin_0128 (RW)
0x6b: frame_modchk_group_bin_0210 (RW)
0x6c: frame_modchk_group_bin_0294 (RW)
0x6d: frame_modchk_group_bin_0052 (RW)
0x6e: frame_modchk_group_bin_0140 (RW)
0x6f: frame_modchk_group_bin_0220 (RW)
0x70: frame_modchk_group_bin_0304 (RW)
0x71: frame_modchk_group_bin_0062 (RW)
0x72: frame_modchk_group_bin_0148 (RW)
0x73: frame_modchk_group_bin_0229 (RW)
0x74: frame_modchk_group_bin_0313 (RW)
0x75: frame_modchk_group_bin_0073 (RW)
0x76: frame_modchk_group_bin_0158 (RW)
0x77: frame_modchk_group_bin_0240 (RW)
0x78: frame_modchk_group_bin_0323 (RW)
0x79: frame_modchk_group_bin_0084 (RW)
0x7: frame_modchk_group_bin_0280 (RX)
0x7a: frame_modchk_group_bin_0168 (RW)
0x7b: frame_modchk_group_bin_0252 (RW)
0x7c: frame_modchk_group_bin_0011 (RW)
0x7d: frame_modchk_group_bin_0095 (RW)
0x7e: frame_modchk_group_bin_0180 (RW)
0x7f: frame_modchk_group_bin_0261 (RW)
0x80: frame_modchk_group_bin_0020 (RW)
0x81: frame_modchk_group_bin_0105 (RW)
0x82: frame_modchk_group_bin_0053 (RW)
0x83: frame_modchk_group_bin_0149 (RW)
0x84: frame_modchk_group_bin_0241 (RW)
0x85: frame_modchk_group_bin_0012 (RW)
0x86: frame_modchk_group_bin_0106 (RW)
0x87: frame_modchk_group_bin_0199 (RW)
0x88: frame_modchk_group_bin_0293 (RW)
0x89: frame_modchk_group_bin_0061 (RW)
0x8: frame_modchk_group_bin_0041 (RX)
0x8a: frame_modchk_group_bin_0157 (RW)
0x8b: frame_modchk_group_bin_0250 (RW)
0x8c: frame_modchk_group_bin_0018 (RW)
0x8d: frame_modchk_group_bin_0117 (RW)
0x8e: frame_modchk_group_bin_0207 (RW)
0x8f: frame_modchk_group_bin_0300 (RW)
0x90: frame_modchk_group_bin_0070 (RW)
0x91: frame_modchk_group_bin_0164 (RW)
0x92: frame_modchk_group_bin_0257 (RW)
0x93: frame_modchk_group_bin_0025 (RW)
0x94: frame_modchk_group_bin_0123 (RW)
0x95: frame_modchk_group_bin_0214 (RW)
0x96: frame_modchk_group_bin_0308 (RW)
0x97: frame_modchk_group_bin_0077 (RW)
0x98: frame_modchk_group_bin_0213 (RW)
0x99: frame_modchk_group_bin_0165 (RW)
0x9: frame_modchk_group_bin_0126 (RX)
0x9a: frame_modchk_group_bin_0181 (RW)
0x9b: frame_modchk_group_bin_0008 (RW)
0x9c: frame_modchk_group_bin_0092 (RW)
0x9d: frame_modchk_group_bin_0286 (RW)
0x9e: frame_modchk_group_bin_0109 (RW)
0x9f: frame_modchk_group_bin_0253 (RW)
0xa0: frame_modchk_group_bin_0273 (RW)
0xa1: frame_modchk_group_bin_0044 (RW)
0xa2: frame_modchk_group_bin_0141 (RW)
0xa3: frame_modchk_group_bin_0230 (RW)
0xa4: frame_modchk_group_bin_0003 (RW)
0xa5: frame_modchk_group_bin_0096 (RW)
0xa6: frame_modchk_group_bin_0190 (RW)
0xa7: frame_modchk_group_bin_0281 (RW)
0xa8: frame_modchk_group_bin_0051 (RW)
0xa9: frame_modchk_group_bin_0147 (RW)
0xa: frame_modchk_group_bin_0208 (RX)
0xaa: frame_modchk_group_bin_0239 (RW)
0xab: frame_modchk_group_bin_0010 (RW)
0xac: frame_modchk_group_bin_0104 (RW)
0xad: frame_modchk_group_bin_0197 (RW)
0xae: frame_modchk_group_bin_0290 (RW)
0xaf: frame_modchk_group_bin_0059 (RW)
0xb0: frame_modchk_group_bin_0154 (RW)
0xb1: frame_modchk_group_bin_0029 (RW)
0xb2: frame_modchk_group_bin_0016 (RW)
0xb3: frame_modchk_group_bin_0114 (RW)
0xb4: frame_modchk_group_bin_0205 (RW)
0xb5: frame_modchk_group_bin_0298 (RW)
0xb6: frame_modchk_group_bin_0067 (RW)
0xb7: frame_modchk_group_bin_0162 (RW)
0xb8: frame_modchk_group_bin_0307 (RW)
0xb9: frame_modchk_group_bin_0129 (RW)
0xb: frame_modchk_group_bin_0291 (RX)
0xba: frame_modchk_group_bin_0005 (RW)
0xbb: frame_modchk_group_bin_0093 (RW)
0xbc: frame_modchk_group_bin_0235 (RW)
0xbd: frame_modchk_group_bin_0056 (RW)
0xbe: frame_modchk_group_bin_0202 (RW)
0xbf: frame_modchk_group_bin_0021 (RW)
0xc0: frame_modchk_group_bin_0032 (RW)
0xc1: frame_modchk_group_bin_0312 (RW)
0xc2: frame_modchk_group_bin_0221 (RW)
0xc3: frame_modchk_group_bin_0314 (RW)
0xc4: frame_modchk_group_bin_0085 (RW)
0xc5: frame_modchk_group_bin_0242 (RW)
0xc6: frame_modchk_group_bin_0271 (RW)
0xc7: frame_modchk_group_bin_0042 (RW)
0xc8: frame_modchk_group_bin_0139 (RW)
0xc9: frame_modchk_group_bin_0228 (RW)
0xc: frame_modchk_group_bin_0049 (RX)
0xca: frame_modchk_group_bin_0322 (RW)
0xcb: frame_modchk_group_bin_0094 (RW)
0xcc: frame_modchk_group_bin_0188 (RW)
0xcd: frame_modchk_group_bin_0279 (RW)
0xce: frame_modchk_group_bin_0048 (RW)
0xcf: frame_modchk_group_bin_0145 (RW)
0xd0: frame_modchk_group_bin_0237 (RW)
0xd1: frame_modchk_group_bin_0007 (RW)
0xd2: frame_modchk_group_bin_0101 (RW)
0xd3: frame_modchk_group_bin_0195 (RW)
0xd4: frame_modchk_group_bin_0288 (RW)
0xd5: frame_modchk_group_bin_0057 (RW)
0xd6: frame_modchk_group_bin_0152 (RW)
0xd7: frame_modchk_group_bin_0245 (RW)
0xd8: frame_modchk_group_bin_0076 (RW)
0xd9: frame_modchk_group_bin_0132 (RW)
0xd: frame_modchk_group_bin_0137 (RX)
0xda: frame_modchk_group_bin_0204 (RW)
0xdb: frame_modchk_group_bin_0187 (RW)
0xdc: frame_modchk_group_bin_0006 (RW)
0xdd: frame_modchk_group_bin_0151 (RW)
0xde: frame_modchk_group_bin_0295 (RW)
0xdf: frame_modchk_group_bin_0119 (RW)
0xe0: frame_modchk_group_bin_0121 (RW)
0xe1: frame_modchk_group_bin_0211 (RW)
0xe2: frame_modchk_group_bin_0305 (RW)
0xe3: frame_modchk_group_bin_0074 (RW)
0xe4: frame_modchk_group_bin_0169 (RW)
0xe5: frame_modchk_group_bin_0262 (RW)
0xe6: frame_modchk_group_bin_0130 (RW)
0xe7: frame_modchk_group_bin_0127 (RW)
0xe8: frame_modchk_group_bin_0218 (RW)
0xe9: frame_modchk_group_bin_0266 (RW)
0xe: frame_modchk_group_bin_0217 (RX)
0xea: frame_modchk_group_bin_0083 (RW)
0xeb: frame_modchk_group_bin_0178 (RW)
0xec: frame_modchk_group_bin_0268 (RW)
0xed: frame_modchk_group_bin_0039 (RW)
0xee: frame_modchk_group_bin_0136 (RW)
0xef: frame_modchk_group_bin_0225 (RW)
0xf0: frame_modchk_group_bin_0320 (RW)
0xf1: frame_modchk_group_bin_0091 (RW)
0xf2: frame_modchk_group_bin_0185 (RW)
0xf3: frame_modchk_group_bin_0276 (RW)
0xf4: frame_modchk_group_bin_0046 (RW)
0xf5: frame_modchk_group_bin_0143 (RW)
0xf6: frame_modchk_group_bin_0233 (RW)
0xf7: frame_modchk_group_bin_0116 (RW)
0xf8: frame_modchk_group_bin_0171 (RW)
0xf9: frame_modchk_group_bin_0274 (RW)
0xf: frame_modchk_group_bin_0301 (RX)
0xfa: frame_modchk_group_bin_0138 (RW)
0xfb: frame_modchk_group_bin_0278 (RW)
0xfc: frame_modchk_group_bin_0100 (RW)
0xfd: frame_modchk_group_bin_0244 (RW)
0xfe: frame_modchk_group_bin_0063 (RW)
0xff: frame_modchk_group_bin_0209 (RW)
}
pt_modtx_group_bin_0002 {
0x0: frame_modtx_group_bin_0000 (RX)
0x100: frame_modtx_group_bin_0030 (RW)
0x101: frame_modtx_group_bin_0178 (RW)
0x102: frame_modtx_group_bin_0231 (RW)
0x103: frame_modtx_group_bin_0159 (RW)
0x104: frame_modtx_group_bin_0283 (RW)
0x105: frame_modtx_group_bin_0107 (RW)
0x106: frame_modtx_group_bin_0250 (RW)
0x107: frame_modtx_group_bin_0296 (RW)
0x108: frame_modtx_group_bin_0302 (RW)
0x109: frame_modtx_group_bin_0072 (RW)
0x10: frame_modtx_group_bin_0060 (RX)
0x10a: frame_modtx_group_bin_0166 (RW)
0x10b: frame_modtx_group_bin_0259 (RW)
0x10c: frame_modtx_group_bin_0027 (RW)
0x10d: frame_modtx_group_bin_0125 (RW)
0x10e: frame_modtx_group_bin_0215 (RW)
0x10f: frame_modtx_group_bin_0309 (RW)
0x110: frame_modtx_group_bin_0080 (RW)
0x111: frame_modtx_group_bin_0175 (RW)
0x112: frame_modtx_group_bin_0111 (RW)
0x113: frame_modtx_group_bin_0037 (RW)
0x114: frame_modtx_group_bin_0133 (RW)
0x115: frame_modtx_group_bin_0222 (RW)
0x116: frame_modtx_group_bin_0317 (RW)
0x117: frame_modtx_group_bin_0089 (RW)
0x118: frame_modtx_group_bin_0263 (RW)
0x119: frame_modtx_group_bin_0086 (RW)
0x11: frame_modtx_group_bin_0146 (RX)
0x11a: frame_modtx_group_bin_0172 (RW)
0x11b: frame_modtx_group_bin_0098 (RW)
0x11c: frame_modtx_group_bin_0193 (RW)
0x11d: frame_modtx_group_bin_0014 (RW)
0x11e: frame_modtx_group_bin_0160 (RW)
0x11f: frame_modtx_group_bin_0190 (RW)
0x120: frame_modtx_group_bin_0282 (RW)
0x121: frame_modtx_group_bin_0268 (RW)
0x122: frame_modtx_group_bin_0235 (RW)
0x123: frame_modtx_group_bin_0024 (RW)
0x124: frame_modtx_group_bin_0054 (RW)
0x125: frame_modtx_group_bin_0199 (RW)
0x126: frame_modtx_group_bin_0019 (RW)
0x127: frame_modtx_group_bin_0291 (RW)
0x129: stack__camkes_stack_modtx_0_control_0_modtx_obj (RW)
0x12: frame_modtx_group_bin_0225 (RX)
0x12a: stack__camkes_stack_modtx_0_control_1_modtx_obj (RW)
0x12b: stack__camkes_stack_modtx_0_control_2_modtx_obj (RW)
0x12c: stack__camkes_stack_modtx_0_control_3_modtx_obj (RW)
0x12f: stack__camkes_stack_modtx_modtx_iface_0000_0_modtx_obj (RW)
0x130: stack__camkes_stack_modtx_modtx_iface_0000_1_modtx_obj (RW)
0x131: stack__camkes_stack_modtx_modtx_iface_0000_2_modtx_obj (RW)
0x132: stack__camkes_stack_modtx_modtx_iface_0000_3_modtx_obj (RW)
0x135: stack__camkes_stack_modtx_0_fault_handler_0000_0_modtx_obj (RW)
0x136: stack__camkes_stack_modtx_0_fault_handler_0000_1_modtx_obj (RW)
0x137: stack__camkes_stack_modtx_0_fault_handler_0000_2_modtx_obj (RW)
0x138: stack__camkes_stack_modtx_0_fault_handler_0000_3_modtx_obj (RW)
0x13: frame_modtx_group_bin_0310 (RX)
0x13b: modtx_frame__camkes_ipc_buffer_modtx_0_control (RW)
0x13e: modtx_frame__camkes_ipc_buffer_modtx_modtx_iface_0000 (RW)
0x141: modtx_frame__camkes_ipc_buffer_modtx_0_fault_handler_0000 (RW)
0x14: frame_modtx_group_bin_0071 (RX)
0x15: frame_modtx_group_bin_0155 (RX)
0x16: frame_modtx_group_bin_0237 (RX)
0x17: frame_modtx_group_bin_0320 (RX)
0x18: frame_modtx_group_bin_0081 (RX)
0x19: frame_modtx_group_bin_0087 (RX)
0x1: frame_modtx_group_bin_0001 (RX)
0x1a: frame_modtx_group_bin_0248 (RX)
0x1b: frame_modtx_group_bin_0247 (RX)
0x1c: frame_modtx_group_bin_0004 (RX)
0x1d: frame_modtx_group_bin_0176 (RX)
0x1e: frame_modtx_group_bin_0257 (RX)
0x1f: frame_modtx_group_bin_0017 (RX)
0x20: frame_modtx_group_bin_0102 (RX)
0x21: frame_modtx_group_bin_0185 (RX)
0x22: frame_modtx_group_bin_0266 (RX)
0x23: frame_modtx_group_bin_0026 (RX)
0x24: frame_modtx_group_bin_0115 (RW)
0x25: frame_modtx_group_bin_0195 (RW)
0x26: frame_modtx_group_bin_0276 (RW)
0x27: frame_modtx_group_bin_0038 (RW)
0x28: frame_modtx_group_bin_0124 (RW)
0x29: frame_modtx_group_bin_0205 (RW)
0x2: frame_modtx_group_bin_0188 (RX)
0x2a: frame_modtx_group_bin_0288 (RW)
0x2b: frame_modtx_group_bin_0047 (RW)
0x2c: frame_modtx_group_bin_0134 (RW)
0x2d: frame_modtx_group_bin_0214 (RW)
0x2e: frame_modtx_group_bin_0298 (RW)
0x2f: frame_modtx_group_bin_0058 (RW)
0x30: frame_modtx_group_bin_0144 (RW)
0x31: frame_modtx_group_bin_0223 (RW)
0x32: frame_modtx_group_bin_0308 (RW)
0x33: frame_modtx_group_bin_0068 (RW)
0x34: frame_modtx_group_bin_0153 (RW)
0x35: frame_modtx_group_bin_0233 (RW)
0x36: frame_modtx_group_bin_0318 (RW)
0x37: frame_modtx_group_bin_0078 (RW)
0x38: frame_modtx_group_bin_0163 (RW)
0x39: frame_modtx_group_bin_0245 (RW)
0x3: frame_modtx_group_bin_0269 (RX)
0x3a: frame_modtx_group_bin_0167 (RW)
0x3b: frame_modtx_group_bin_0090 (RW)
0x3c: frame_modtx_group_bin_0173 (RW)
0x3d: frame_modtx_group_bin_0255 (RW)
0x3e: frame_modtx_group_bin_0015 (RW)
0x3f: frame_modtx_group_bin_0099 (RW)
0x40: frame_modtx_group_bin_0183 (RW)
0x41: frame_modtx_group_bin_0264 (RW)
0x42: frame_modtx_group_bin_0023 (RW)
0x43: frame_modtx_group_bin_0112 (RW)
0x44: frame_modtx_group_bin_0192 (RW)
0x45: frame_modtx_group_bin_0274 (RW)
0x46: frame_modtx_group_bin_0035 (RW)
0x47: frame_modtx_group_bin_0122 (RW)
0x48: frame_modtx_group_bin_0202 (RW)
0x49: frame_modtx_group_bin_0284 (RW)
0x4: frame_modtx_group_bin_0028 (RX)
0x4a: frame_modtx_group_bin_0045 (RW)
0x4b: frame_modtx_group_bin_0131 (RW)
0x4c: frame_modtx_group_bin_0211 (RW)
0x4d: frame_modtx_group_bin_0295 (RW)
0x4e: frame_modtx_group_bin_0055 (RW)
0x4f: frame_modtx_group_bin_0142 (RW)
0x50: frame_modtx_group_bin_0221 (RW)
0x51: frame_modtx_group_bin_0305 (RW)
0x52: frame_modtx_group_bin_0065 (RW)
0x53: frame_modtx_group_bin_0150 (RW)
0x54: frame_modtx_group_bin_0230 (RW)
0x55: frame_modtx_group_bin_0315 (RW)
0x56: frame_modtx_group_bin_0075 (RW)
0x57: frame_modtx_group_bin_0161 (RW)
0x58: frame_modtx_group_bin_0242 (RW)
0x59: frame_modtx_group_bin_0002 (RW)
0x5: frame_modtx_group_bin_0118 (RX)
0x5a: frame_modtx_group_bin_0088 (RW)
0x5b: frame_modtx_group_bin_0170 (RW)
0x5c: frame_modtx_group_bin_0254 (RW)
0x5d: frame_modtx_group_bin_0013 (RW)
0x5e: frame_modtx_group_bin_0097 (RW)
0x5f: frame_modtx_group_bin_0182 (RW)
0x60: frame_modtx_group_bin_0262 (RW)
0x61: frame_modtx_group_bin_0022 (RW)
0x62: frame_modtx_group_bin_0108 (RW)
0x63: frame_modtx_group_bin_0191 (RW)
0x64: frame_modtx_group_bin_0271 (RW)
0x65: frame_modtx_group_bin_0031 (RW)
0x66: frame_modtx_group_bin_0120 (RW)
0x67: frame_modtx_group_bin_0200 (RW)
0x68: frame_modtx_group_bin_0281 (RW)
0x69: frame_modtx_group_bin_0043 (RW)
0x6: frame_modtx_group_bin_0197 (RX)
0x6a: frame_modtx_group_bin_0128 (RW)
0x6b: frame_modtx_group_bin_0209 (RW)
0x6c: frame_modtx_group_bin_0293 (RW)
0x6d: frame_modtx_group_bin_0052 (RW)
0x6e: frame_modtx_group_bin_0140 (RW)
0x6f: frame_modtx_group_bin_0219 (RW)
0x70: frame_modtx_group_bin_0303 (RW)
0x71: frame_modtx_group_bin_0062 (RW)
0x72: frame_modtx_group_bin_0148 (RW)
0x73: frame_modtx_group_bin_0228 (RW)
0x74: frame_modtx_group_bin_0312 (RW)
0x75: frame_modtx_group_bin_0073 (RW)
0x76: frame_modtx_group_bin_0158 (RW)
0x77: frame_modtx_group_bin_0239 (RW)
0x78: frame_modtx_group_bin_0322 (RW)
0x79: frame_modtx_group_bin_0084 (RW)
0x7: frame_modtx_group_bin_0279 (RX)
0x7a: frame_modtx_group_bin_0168 (RW)
0x7b: frame_modtx_group_bin_0251 (RW)
0x7c: frame_modtx_group_bin_0011 (RW)
0x7d: frame_modtx_group_bin_0095 (RW)
0x7e: frame_modtx_group_bin_0179 (RW)
0x7f: frame_modtx_group_bin_0260 (RW)
0x80: frame_modtx_group_bin_0020 (RW)
0x81: frame_modtx_group_bin_0105 (RW)
0x82: frame_modtx_group_bin_0053 (RW)
0x83: frame_modtx_group_bin_0149 (RW)
0x84: frame_modtx_group_bin_0240 (RW)
0x85: frame_modtx_group_bin_0012 (RW)
0x86: frame_modtx_group_bin_0106 (RW)
0x87: frame_modtx_group_bin_0198 (RW)
0x88: frame_modtx_group_bin_0292 (RW)
0x89: frame_modtx_group_bin_0061 (RW)
0x8: frame_modtx_group_bin_0041 (RX)
0x8a: frame_modtx_group_bin_0157 (RW)
0x8b: frame_modtx_group_bin_0249 (RW)
0x8c: frame_modtx_group_bin_0018 (RW)
0x8d: frame_modtx_group_bin_0117 (RW)
0x8e: frame_modtx_group_bin_0206 (RW)
0x8f: frame_modtx_group_bin_0299 (RW)
0x90: frame_modtx_group_bin_0070 (RW)
0x91: frame_modtx_group_bin_0164 (RW)
0x92: frame_modtx_group_bin_0256 (RW)
0x93: frame_modtx_group_bin_0025 (RW)
0x94: frame_modtx_group_bin_0123 (RW)
0x95: frame_modtx_group_bin_0213 (RW)
0x96: frame_modtx_group_bin_0307 (RW)
0x97: frame_modtx_group_bin_0077 (RW)
0x98: frame_modtx_group_bin_0212 (RW)
0x99: frame_modtx_group_bin_0165 (RW)
0x9: frame_modtx_group_bin_0126 (RX)
0x9a: frame_modtx_group_bin_0180 (RW)
0x9b: frame_modtx_group_bin_0008 (RW)
0x9c: frame_modtx_group_bin_0092 (RW)
0x9d: frame_modtx_group_bin_0285 (RW)
0x9e: frame_modtx_group_bin_0109 (RW)
0x9f: frame_modtx_group_bin_0252 (RW)
0xa0: frame_modtx_group_bin_0272 (RW)
0xa1: frame_modtx_group_bin_0044 (RW)
0xa2: frame_modtx_group_bin_0141 (RW)
0xa3: frame_modtx_group_bin_0229 (RW)
0xa4: frame_modtx_group_bin_0003 (RW)
0xa5: frame_modtx_group_bin_0096 (RW)
0xa6: frame_modtx_group_bin_0189 (RW)
0xa7: frame_modtx_group_bin_0280 (RW)
0xa8: frame_modtx_group_bin_0051 (RW)
0xa9: frame_modtx_group_bin_0147 (RW)
0xa: frame_modtx_group_bin_0207 (RX)
0xaa: frame_modtx_group_bin_0238 (RW)
0xab: frame_modtx_group_bin_0010 (RW)
0xac: frame_modtx_group_bin_0104 (RW)
0xad: frame_modtx_group_bin_0196 (RW)
0xae: frame_modtx_group_bin_0289 (RW)
0xaf: frame_modtx_group_bin_0059 (RW)
0xb0: frame_modtx_group_bin_0154 (RW)
0xb1: frame_modtx_group_bin_0029 (RW)
0xb2: frame_modtx_group_bin_0016 (RW)
0xb3: frame_modtx_group_bin_0114 (RW)
0xb4: frame_modtx_group_bin_0204 (RW)
0xb5: frame_modtx_group_bin_0297 (RW)
0xb6: frame_modtx_group_bin_0067 (RW)
0xb7: frame_modtx_group_bin_0162 (RW)
0xb8: frame_modtx_group_bin_0306 (RW)
0xb9: frame_modtx_group_bin_0129 (RW)
0xb: frame_modtx_group_bin_0290 (RX)
0xba: frame_modtx_group_bin_0005 (RW)
0xbb: frame_modtx_group_bin_0093 (RW)
0xbc: frame_modtx_group_bin_0234 (RW)
0xbd: frame_modtx_group_bin_0056 (RW)
0xbe: frame_modtx_group_bin_0201 (RW)
0xbf: frame_modtx_group_bin_0021 (RW)
0xc0: frame_modtx_group_bin_0032 (RW)
0xc1: frame_modtx_group_bin_0311 (RW)
0xc2: frame_modtx_group_bin_0220 (RW)
0xc3: frame_modtx_group_bin_0313 (RW)
0xc4: frame_modtx_group_bin_0085 (RW)
0xc5: frame_modtx_group_bin_0241 (RW)
0xc6: frame_modtx_group_bin_0270 (RW)
0xc7: frame_modtx_group_bin_0042 (RW)
0xc8: frame_modtx_group_bin_0139 (RW)
0xc9: frame_modtx_group_bin_0227 (RW)
0xc: frame_modtx_group_bin_0049 (RX)
0xca: frame_modtx_group_bin_0321 (RW)
0xcb: frame_modtx_group_bin_0094 (RW)
0xcc: frame_modtx_group_bin_0187 (RW)
0xcd: frame_modtx_group_bin_0278 (RW)
0xce: frame_modtx_group_bin_0048 (RW)
0xcf: frame_modtx_group_bin_0145 (RW)
0xd0: frame_modtx_group_bin_0236 (RW)
0xd1: frame_modtx_group_bin_0007 (RW)
0xd2: frame_modtx_group_bin_0101 (RW)
0xd3: frame_modtx_group_bin_0194 (RW)
0xd4: frame_modtx_group_bin_0287 (RW)
0xd5: frame_modtx_group_bin_0057 (RW)
0xd6: frame_modtx_group_bin_0152 (RW)
0xd7: frame_modtx_group_bin_0244 (RW)
0xd8: frame_modtx_group_bin_0076 (RW)
0xd9: frame_modtx_group_bin_0132 (RW)
0xd: frame_modtx_group_bin_0137 (RX)
0xda: frame_modtx_group_bin_0203 (RW)
0xdb: frame_modtx_group_bin_0186 (RW)
0xdc: frame_modtx_group_bin_0006 (RW)
0xdd: frame_modtx_group_bin_0151 (RW)
0xde: frame_modtx_group_bin_0294 (RW)
0xdf: frame_modtx_group_bin_0119 (RW)
0xe0: frame_modtx_group_bin_0121 (RW)
0xe1: frame_modtx_group_bin_0210 (RW)
0xe2: frame_modtx_group_bin_0304 (RW)
0xe3: frame_modtx_group_bin_0074 (RW)
0xe4: frame_modtx_group_bin_0169 (RW)
0xe5: frame_modtx_group_bin_0261 (RW)
0xe6: frame_modtx_group_bin_0130 (RW)
0xe7: frame_modtx_group_bin_0127 (RW)
0xe8: frame_modtx_group_bin_0217 (RW)
0xe9: frame_modtx_group_bin_0265 (RW)
0xe: frame_modtx_group_bin_0216 (RX)
0xea: frame_modtx_group_bin_0083 (RW)
0xeb: frame_modtx_group_bin_0177 (RW)
0xec: frame_modtx_group_bin_0267 (RW)
0xed: frame_modtx_group_bin_0039 (RW)
0xee: frame_modtx_group_bin_0136 (RW)
0xef: frame_modtx_group_bin_0224 (RW)
0xf0: frame_modtx_group_bin_0319 (RW)
0xf1: frame_modtx_group_bin_0091 (RW)
0xf2: frame_modtx_group_bin_0184 (RW)
0xf3: frame_modtx_group_bin_0275 (RW)
0xf4: frame_modtx_group_bin_0046 (RW)
0xf5: frame_modtx_group_bin_0143 (RW)
0xf6: frame_modtx_group_bin_0232 (RW)
0xf7: frame_modtx_group_bin_0116 (RW)
0xf8: frame_modtx_group_bin_0171 (RW)
0xf9: frame_modtx_group_bin_0273 (RW)
0xf: frame_modtx_group_bin_0300 (RX)
0xfa: frame_modtx_group_bin_0138 (RW)
0xfb: frame_modtx_group_bin_0277 (RW)
0xfc: frame_modtx_group_bin_0100 (RW)
0xfd: frame_modtx_group_bin_0243 (RW)
0xfe: frame_modtx_group_bin_0063 (RW)
0xff: frame_modtx_group_bin_0208 (RW)
}
pt_signtx_group_bin_0002 {
0x0: frame_signtx_group_bin_0000 (RX)
0x100: frame_signtx_group_bin_0030 (RW)
0x101: frame_signtx_group_bin_0180 (RW)
0x102: frame_signtx_group_bin_0233 (RW)
0x103: frame_signtx_group_bin_0160 (RW)
0x104: frame_signtx_group_bin_0285 (RW)
0x105: frame_signtx_group_bin_0107 (RW)
0x106: frame_signtx_group_bin_0252 (RW)
0x107: frame_signtx_group_bin_0298 (RW)
0x108: frame_signtx_group_bin_0304 (RW)
0x109: frame_signtx_group_bin_0072 (RW)
0x10: frame_signtx_group_bin_0060 (RX)
0x10a: frame_signtx_group_bin_0167 (RW)
0x10b: frame_signtx_group_bin_0261 (RW)
0x10c: frame_signtx_group_bin_0027 (RW)
0x10d: frame_signtx_group_bin_0125 (RW)
0x10e: frame_signtx_group_bin_0217 (RW)
0x10f: frame_signtx_group_bin_0311 (RW)
0x110: frame_signtx_group_bin_0080 (RW)
0x111: frame_signtx_group_bin_0177 (RW)
0x112: frame_signtx_group_bin_0111 (RW)
0x113: frame_signtx_group_bin_0037 (RW)
0x114: frame_signtx_group_bin_0133 (RW)
0x115: frame_signtx_group_bin_0224 (RW)
0x116: frame_signtx_group_bin_0319 (RW)
0x117: frame_signtx_group_bin_0089 (RW)
0x118: frame_signtx_group_bin_0265 (RW)
0x119: frame_signtx_group_bin_0086 (RW)
0x11: frame_signtx_group_bin_0146 (RX)
0x11a: frame_signtx_group_bin_0174 (RW)
0x11b: frame_signtx_group_bin_0098 (RW)
0x11c: frame_signtx_group_bin_0195 (RW)
0x11d: frame_signtx_group_bin_0014 (RW)
0x11e: frame_signtx_group_bin_0161 (RW)
0x11f: frame_signtx_group_bin_0192 (RW)
0x120: frame_signtx_group_bin_0284 (RW)
0x121: frame_signtx_group_bin_0270 (RW)
0x122: frame_signtx_group_bin_0237 (RW)
0x123: frame_signtx_group_bin_0024 (RW)
0x124: frame_signtx_group_bin_0054 (RW)
0x125: frame_signtx_group_bin_0201 (RW)
0x126: frame_signtx_group_bin_0019 (RW)
0x127: frame_signtx_group_bin_0293 (RW)
0x128: frame_signtx_group_bin_0260 (RW)
0x129: frame_signtx_group_bin_0009 (RW)
0x12: frame_signtx_group_bin_0227 (RX)
0x12b: stack__camkes_stack_signtx_0_control_0_signtx_obj (RW)
0x12c: stack__camkes_stack_signtx_0_control_1_signtx_obj (RW)
0x12d: stack__camkes_stack_signtx_0_control_2_signtx_obj (RW)
0x12e: stack__camkes_stack_signtx_0_control_3_signtx_obj (RW)
0x131: stack__camkes_stack_signtx_signtx_iface_0000_0_signtx_obj (RW)
0x132: stack__camkes_stack_signtx_signtx_iface_0000_1_signtx_obj (RW)
0x133: stack__camkes_stack_signtx_signtx_iface_0000_2_signtx_obj (RW)
0x134: stack__camkes_stack_signtx_signtx_iface_0000_3_signtx_obj (RW)
0x137: stack__camkes_stack_signtx_0_fault_handler_0000_0_signtx_obj (RW)
0x138: stack__camkes_stack_signtx_0_fault_handler_0000_1_signtx_obj (RW)
0x139: stack__camkes_stack_signtx_0_fault_handler_0000_2_signtx_obj (RW)
0x13: frame_signtx_group_bin_0312 (RX)
0x13a: stack__camkes_stack_signtx_0_fault_handler_0000_3_signtx_obj (RW)
0x13d: signtx_frame__camkes_ipc_buffer_signtx_0_control (RW)
0x140: signtx_frame__camkes_ipc_buffer_signtx_signtx_iface_0000 (RW)
0x143: signtx_frame__camkes_ipc_buffer_signtx_0_fault_handler_0000 (RW)
0x14: frame_signtx_group_bin_0071 (RX)
0x15: frame_signtx_group_bin_0156 (RX)
0x16: frame_signtx_group_bin_0239 (RX)
0x17: frame_signtx_group_bin_0322 (RX)
0x18: frame_signtx_group_bin_0081 (RX)
0x19: frame_signtx_group_bin_0087 (RX)
0x1: frame_signtx_group_bin_0001 (RX)
0x1a: frame_signtx_group_bin_0250 (RX)
0x1b: frame_signtx_group_bin_0249 (RX)
0x1c: frame_signtx_group_bin_0004 (RX)
0x1d: frame_signtx_group_bin_0178 (RX)
0x1e: frame_signtx_group_bin_0259 (RX)
0x1f: frame_signtx_group_bin_0017 (RX)
0x20: frame_signtx_group_bin_0102 (RX)
0x21: frame_signtx_group_bin_0187 (RX)
0x22: frame_signtx_group_bin_0268 (RX)
0x23: frame_signtx_group_bin_0026 (RX)
0x24: frame_signtx_group_bin_0115 (RX)
0x25: frame_signtx_group_bin_0197 (RX)
0x26: frame_signtx_group_bin_0278 (RW)
0x27: frame_signtx_group_bin_0038 (RW)
0x28: frame_signtx_group_bin_0124 (RW)
0x29: frame_signtx_group_bin_0207 (RW)
0x2: frame_signtx_group_bin_0190 (RX)
0x2a: frame_signtx_group_bin_0290 (RW)
0x2b: frame_signtx_group_bin_0047 (RW)
0x2c: frame_signtx_group_bin_0134 (RW)
0x2d: frame_signtx_group_bin_0216 (RW)
0x2e: frame_signtx_group_bin_0300 (RW)
0x2f: frame_signtx_group_bin_0058 (RW)
0x30: frame_signtx_group_bin_0144 (RW)
0x31: frame_signtx_group_bin_0225 (RW)
0x32: frame_signtx_group_bin_0310 (RW)
0x33: frame_signtx_group_bin_0068 (RW)
0x34: frame_signtx_group_bin_0154 (RW)
0x35: frame_signtx_group_bin_0235 (RW)
0x36: frame_signtx_group_bin_0320 (RW)
0x37: frame_signtx_group_bin_0078 (RW)
0x38: frame_signtx_group_bin_0164 (RW)
0x39: frame_signtx_group_bin_0247 (RW)
0x3: frame_signtx_group_bin_0271 (RX)
0x3a: frame_signtx_group_bin_0168 (RW)
0x3b: frame_signtx_group_bin_0090 (RW)
0x3c: frame_signtx_group_bin_0175 (RW)
0x3d: frame_signtx_group_bin_0257 (RW)
0x3e: frame_signtx_group_bin_0015 (RW)
0x3f: frame_signtx_group_bin_0099 (RW)
0x40: frame_signtx_group_bin_0185 (RW)
0x41: frame_signtx_group_bin_0266 (RW)
0x42: frame_signtx_group_bin_0023 (RW)
0x43: frame_signtx_group_bin_0112 (RW)
0x44: frame_signtx_group_bin_0194 (RW)
0x45: frame_signtx_group_bin_0276 (RW)
0x46: frame_signtx_group_bin_0035 (RW)
0x47: frame_signtx_group_bin_0122 (RW)
0x48: frame_signtx_group_bin_0204 (RW)
0x49: frame_signtx_group_bin_0286 (RW)
0x4: frame_signtx_group_bin_0028 (RX)
0x4a: frame_signtx_group_bin_0045 (RW)
0x4b: frame_signtx_group_bin_0131 (RW)
0x4c: frame_signtx_group_bin_0213 (RW)
0x4d: frame_signtx_group_bin_0297 (RW)
0x4e: frame_signtx_group_bin_0055 (RW)
0x4f: frame_signtx_group_bin_0142 (RW)
0x50: frame_signtx_group_bin_0223 (RW)
0x51: frame_signtx_group_bin_0307 (RW)
0x52: frame_signtx_group_bin_0065 (RW)
0x53: frame_signtx_group_bin_0151 (RW)
0x54: frame_signtx_group_bin_0232 (RW)
0x55: frame_signtx_group_bin_0317 (RW)
0x56: frame_signtx_group_bin_0075 (RW)
0x57: frame_signtx_group_bin_0162 (RW)
0x58: frame_signtx_group_bin_0244 (RW)
0x59: frame_signtx_group_bin_0002 (RW)
0x5: frame_signtx_group_bin_0118 (RX)
0x5a: frame_signtx_group_bin_0088 (RW)
0x5b: frame_signtx_group_bin_0171 (RW)
0x5c: frame_signtx_group_bin_0256 (RW)
0x5d: frame_signtx_group_bin_0013 (RW)
0x5e: frame_signtx_group_bin_0097 (RW)
0x5f: frame_signtx_group_bin_0184 (RW)
0x60: frame_signtx_group_bin_0264 (RW)
0x61: frame_signtx_group_bin_0022 (RW)
0x62: frame_signtx_group_bin_0108 (RW)
0x63: frame_signtx_group_bin_0193 (RW)
0x64: frame_signtx_group_bin_0273 (RW)
0x65: frame_signtx_group_bin_0031 (RW)
0x66: frame_signtx_group_bin_0120 (RW)
0x67: frame_signtx_group_bin_0202 (RW)
0x68: frame_signtx_group_bin_0283 (RW)
0x69: frame_signtx_group_bin_0043 (RW)
0x6: frame_signtx_group_bin_0199 (RX)
0x6a: frame_signtx_group_bin_0128 (RW)
0x6b: frame_signtx_group_bin_0211 (RW)
0x6c: frame_signtx_group_bin_0295 (RW)
0x6d: frame_signtx_group_bin_0052 (RW)
0x6e: frame_signtx_group_bin_0140 (RW)
0x6f: frame_signtx_group_bin_0221 (RW)
0x70: frame_signtx_group_bin_0305 (RW)
0x71: frame_signtx_group_bin_0062 (RW)
0x72: frame_signtx_group_bin_0148 (RW)
0x73: frame_signtx_group_bin_0230 (RW)
0x74: frame_signtx_group_bin_0314 (RW)
0x75: frame_signtx_group_bin_0073 (RW)
0x76: frame_signtx_group_bin_0159 (RW)
0x77: frame_signtx_group_bin_0241 (RW)
0x78: frame_signtx_group_bin_0324 (RW)
0x79: frame_signtx_group_bin_0084 (RW)
0x7: frame_signtx_group_bin_0281 (RX)
0x7a: frame_signtx_group_bin_0169 (RW)
0x7b: frame_signtx_group_bin_0253 (RW)
0x7c: frame_signtx_group_bin_0011 (RW)
0x7d: frame_signtx_group_bin_0095 (RW)
0x7e: frame_signtx_group_bin_0181 (RW)
0x7f: frame_signtx_group_bin_0262 (RW)
0x80: frame_signtx_group_bin_0020 (RW)
0x81: frame_signtx_group_bin_0105 (RW)
0x82: frame_signtx_group_bin_0053 (RW)
0x83: frame_signtx_group_bin_0149 (RW)
0x84: frame_signtx_group_bin_0242 (RW)
0x85: frame_signtx_group_bin_0012 (RW)
0x86: frame_signtx_group_bin_0106 (RW)
0x87: frame_signtx_group_bin_0200 (RW)
0x88: frame_signtx_group_bin_0294 (RW)
0x89: frame_signtx_group_bin_0061 (RW)
0x8: frame_signtx_group_bin_0041 (RX)
0x8a: frame_signtx_group_bin_0158 (RW)
0x8b: frame_signtx_group_bin_0251 (RW)
0x8c: frame_signtx_group_bin_0018 (RW)
0x8d: frame_signtx_group_bin_0117 (RW)
0x8e: frame_signtx_group_bin_0208 (RW)
0x8f: frame_signtx_group_bin_0301 (RW)
0x90: frame_signtx_group_bin_0070 (RW)
0x91: frame_signtx_group_bin_0165 (RW)
0x92: frame_signtx_group_bin_0258 (RW)
0x93: frame_signtx_group_bin_0025 (RW)
0x94: frame_signtx_group_bin_0123 (RW)
0x95: frame_signtx_group_bin_0215 (RW)
0x96: frame_signtx_group_bin_0309 (RW)
0x97: frame_signtx_group_bin_0077 (RW)
0x98: frame_signtx_group_bin_0214 (RW)
0x99: frame_signtx_group_bin_0166 (RW)
0x9: frame_signtx_group_bin_0126 (RX)
0x9a: frame_signtx_group_bin_0182 (RW)
0x9b: frame_signtx_group_bin_0008 (RW)
0x9c: frame_signtx_group_bin_0092 (RW)
0x9d: frame_signtx_group_bin_0287 (RW)
0x9e: frame_signtx_group_bin_0109 (RW)
0x9f: frame_signtx_group_bin_0254 (RW)
0xa0: frame_signtx_group_bin_0274 (RW)
0xa1: frame_signtx_group_bin_0044 (RW)
0xa2: frame_signtx_group_bin_0141 (RW)
0xa3: frame_signtx_group_bin_0231 (RW)
0xa4: frame_signtx_group_bin_0003 (RW)
0xa5: frame_signtx_group_bin_0096 (RW)
0xa6: frame_signtx_group_bin_0191 (RW)
0xa7: frame_signtx_group_bin_0282 (RW)
0xa8: frame_signtx_group_bin_0051 (RW)
0xa9: frame_signtx_group_bin_0147 (RW)
0xa: frame_signtx_group_bin_0209 (RX)
0xaa: frame_signtx_group_bin_0240 (RW)
0xab: frame_signtx_group_bin_0010 (RW)
0xac: frame_signtx_group_bin_0104 (RW)
0xad: frame_signtx_group_bin_0198 (RW)
0xae: frame_signtx_group_bin_0291 (RW)
0xaf: frame_signtx_group_bin_0059 (RW)
0xb0: frame_signtx_group_bin_0155 (RW)
0xb1: frame_signtx_group_bin_0029 (RW)
0xb2: frame_signtx_group_bin_0016 (RW)
0xb3: frame_signtx_group_bin_0114 (RW)
0xb4: frame_signtx_group_bin_0206 (RW)
0xb5: frame_signtx_group_bin_0299 (RW)
0xb6: frame_signtx_group_bin_0067 (RW)
0xb7: frame_signtx_group_bin_0163 (RW)
0xb8: frame_signtx_group_bin_0308 (RW)
0xb9: frame_signtx_group_bin_0129 (RW)
0xb: frame_signtx_group_bin_0292 (RX)
0xba: frame_signtx_group_bin_0005 (RW)
0xbb: frame_signtx_group_bin_0093 (RW)
0xbc: frame_signtx_group_bin_0236 (RW)
0xbd: frame_signtx_group_bin_0056 (RW)
0xbe: frame_signtx_group_bin_0203 (RW)
0xbf: frame_signtx_group_bin_0021 (RW)
0xc0: frame_signtx_group_bin_0032 (RW)
0xc1: frame_signtx_group_bin_0313 (RW)
0xc2: frame_signtx_group_bin_0222 (RW)
0xc3: frame_signtx_group_bin_0315 (RW)
0xc4: frame_signtx_group_bin_0085 (RW)
0xc5: frame_signtx_group_bin_0243 (RW)
0xc6: frame_signtx_group_bin_0272 (RW)
0xc7: frame_signtx_group_bin_0042 (RW)
0xc8: frame_signtx_group_bin_0139 (RW)
0xc9: frame_signtx_group_bin_0229 (RW)
0xc: frame_signtx_group_bin_0049 (RX)
0xca: frame_signtx_group_bin_0323 (RW)
0xcb: frame_signtx_group_bin_0094 (RW)
0xcc: frame_signtx_group_bin_0189 (RW)
0xcd: frame_signtx_group_bin_0280 (RW)
0xce: frame_signtx_group_bin_0048 (RW)
0xcf: frame_signtx_group_bin_0145 (RW)
0xd0: frame_signtx_group_bin_0238 (RW)
0xd1: frame_signtx_group_bin_0007 (RW)
0xd2: frame_signtx_group_bin_0101 (RW)
0xd3: frame_signtx_group_bin_0196 (RW)
0xd4: frame_signtx_group_bin_0289 (RW)
0xd5: frame_signtx_group_bin_0057 (RW)
0xd6: frame_signtx_group_bin_0153 (RW)
0xd7: frame_signtx_group_bin_0246 (RW)
0xd8: frame_signtx_group_bin_0076 (RW)
0xd9: frame_signtx_group_bin_0132 (RW)
0xd: frame_signtx_group_bin_0137 (RX)
0xda: frame_signtx_group_bin_0205 (RW)
0xdb: frame_signtx_group_bin_0188 (RW)
0xdc: frame_signtx_group_bin_0006 (RW)
0xdd: frame_signtx_group_bin_0152 (RW)
0xde: frame_signtx_group_bin_0296 (RW)
0xdf: frame_signtx_group_bin_0119 (RW)
0xe0: frame_signtx_group_bin_0121 (RW)
0xe1: frame_signtx_group_bin_0212 (RW)
0xe2: frame_signtx_group_bin_0306 (RW)
0xe3: frame_signtx_group_bin_0074 (RW)
0xe4: frame_signtx_group_bin_0170 (RW)
0xe5: frame_signtx_group_bin_0263 (RW)
0xe6: frame_signtx_group_bin_0130 (RW)
0xe7: frame_signtx_group_bin_0127 (RW)
0xe8: frame_signtx_group_bin_0219 (RW)
0xe9: frame_signtx_group_bin_0267 (RW)
0xe: frame_signtx_group_bin_0218 (RX)
0xea: frame_signtx_group_bin_0083 (RW)
0xeb: frame_signtx_group_bin_0179 (RW)
0xec: frame_signtx_group_bin_0269 (RW)
0xed: frame_signtx_group_bin_0039 (RW)
0xee: frame_signtx_group_bin_0136 (RW)
0xef: frame_signtx_group_bin_0226 (RW)
0xf0: frame_signtx_group_bin_0321 (RW)
0xf1: frame_signtx_group_bin_0091 (RW)
0xf2: frame_signtx_group_bin_0186 (RW)
0xf3: frame_signtx_group_bin_0277 (RW)
0xf4: frame_signtx_group_bin_0046 (RW)
0xf5: frame_signtx_group_bin_0143 (RW)
0xf6: frame_signtx_group_bin_0234 (RW)
0xf7: frame_signtx_group_bin_0116 (RW)
0xf8: frame_signtx_group_bin_0172 (RW)
0xf9: frame_signtx_group_bin_0275 (RW)
0xf: frame_signtx_group_bin_0302 (RX)
0xfa: frame_signtx_group_bin_0138 (RW)
0xfb: frame_signtx_group_bin_0279 (RW)
0xfc: frame_signtx_group_bin_0100 (RW)
0xfd: frame_signtx_group_bin_0245 (RW)
0xfe: frame_signtx_group_bin_0063 (RW)
0xff: frame_signtx_group_bin_0210 (RW)
}
signtx_6_0_control_9_tcb {
cspace: signtx_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: signtx_frame__camkes_ipc_buffer_signtx_0_control (RW)
vspace: signtx_group_bin_pd
}
signtx_6_0_fault_handler_15_0000_tcb {
cspace: signtx_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: signtx_frame__camkes_ipc_buffer_signtx_0_fault_handler_0000 (RW)
vspace: signtx_group_bin_pd
}
signtx_6_signtx_iface_12_0000_tcb {
cspace: signtx_cnode (guard: 0, guard_size: 60)
ipc_buffer_slot: signtx_frame__camkes_ipc_buffer_signtx_signtx_iface_0000 (RW)
vspace: signtx_group_bin_pd
}
signtx_cnode {
0x1: signtx_6_0_control_9_tcb
0x2: signtx_fault_ep (RWX, badge: 1)
0x3: signtx_6_signtx_iface_12_0000_tcb
0x4: signtx_fault_ep (RWX, badge: 3)
0x5: signtx_6_0_fault_handler_15_0000_tcb
0x6: signtx_fault_ep (RWX)
0x7: signtx_pre_init_ep (RW)
0x8: signtx_interface_init_ep (RW)
0x9: signtx_post_init_ep (RW)
0xa: conn2.conn5_ep (WX, badge: 2)
0xb: conn1.conn6_ep (WX, badge: 2)
0xc: conn4.conn8_ep (RW)
0xd: signtx_cnode (guard: 0, guard_size: 60)
}
signtx_group_bin_pd {
0x0: pdpt_signtx_group_bin_0000
}
}

irq maps {

}